* NGSPICE file created from tempsenseInst_error.ext - technology: sky130A

.subckt HEADER VIN sky130_fd_sc_hd__tap_1_1/VPB a_508_138# VGND VNB VPWR sky130_fd_sc_hd__tap_1_0/VPB
X0 a_508_138# VGND VPWR VNB sky130_fd_pr__nfet_03v3_nvt ad=1.1445e+12p pd=1.167e+07u as=3.92e+11p ps=3.92e+06u w=700000u l=500000u
X1 VIN VGND a_508_138# VNB sky130_fd_pr__nfet_03v3_nvt ad=3.92e+11p pd=3.92e+06u as=0p ps=0u w=700000u l=500000u
X2 VPWR VGND a_508_138# VNB sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X3 a_508_138# VGND VPWR VNB sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X4 a_508_138# VGND VIN VNB sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X5 VPWR VGND a_508_138# VNB sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X6 a_508_138# VGND VIN VNB sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
X7 VIN VGND a_508_138# VNB sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=700000u l=500000u
C0 a_508_138# VPWR 0.18fF
C1 a_508_138# VGND 0.56fF
C2 sky130_fd_sc_hd__tap_1_1/VPB VIN 0.00fF
C3 VGND VPWR 0.56fF
C4 VIN sky130_fd_sc_hd__tap_1_0/VPB 0.00fF
C5 sky130_fd_sc_hd__tap_1_1/VPB a_508_138# 0.00fF
C6 a_508_138# sky130_fd_sc_hd__tap_1_0/VPB 0.00fF
C7 sky130_fd_sc_hd__tap_1_1/VPB VPWR 0.07fF
C8 sky130_fd_sc_hd__tap_1_1/VPB VGND 0.02fF
C9 a_508_138# VIN 0.28fF
C10 VPWR sky130_fd_sc_hd__tap_1_0/VPB 0.05fF
C11 VGND sky130_fd_sc_hd__tap_1_0/VPB 0.04fF
C12 VPWR VIN 0.21fF
C13 VGND VIN 0.67fF
C14 VIN VNB 0.61fF
C15 a_508_138# VNB 0.11fF
C16 sky130_fd_sc_hd__tap_1_0/VPB VNB 0.32fF
C17 VGND VNB 3.17fF
C18 VPWR VNB 1.59fF
C19 sky130_fd_sc_hd__tap_1_1/VPB VNB 0.31fF
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=1.05e+06u
C0 VPWR VPB 0.07fF
C1 VPB VGND 0.05fF
C2 VPWR VGND 0.52fF
C3 VPWR VNB 0.61fF
C4 VGND VNB 0.56fF
C5 VPB VNB 0.43fF
.ends

.subckt sky130_fd_sc_hd__or3_1 A X B C VPWR VGND a_29_53# a_183_297# VNB VPB a_111_297#
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=2.965e+11p ps=2.68e+06u w=1e+06u l=150000u
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=3.1715e+11p ps=3.36e+06u w=650000u l=150000u
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=2.226e+11p pd=2.74e+06u as=0p ps=0u w=420000u l=150000u
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 VGND C 0.01fF
C1 a_29_53# B 0.10fF
C2 VPWR a_29_53# 0.07fF
C3 VGND B 0.01fF
C4 a_183_297# A 0.00fF
C5 VGND VPWR 0.05fF
C6 C B 0.06fF
C7 C VPWR 0.00fF
C8 a_183_297# a_29_53# 0.00fF
C9 VGND a_183_297# 0.00fF
C10 VPWR B 0.11fF
C11 a_111_297# A 0.00fF
C12 a_29_53# a_111_297# 0.00fF
C13 X VPB 0.01fF
C14 a_183_297# B 0.00fF
C15 VGND a_111_297# 0.00fF
C16 VPWR a_183_297# 0.00fF
C17 B a_111_297# 0.00fF
C18 VPWR a_111_297# 0.00fF
C19 X A 0.00fF
C20 X a_29_53# 0.07fF
C21 VPB A 0.01fF
C22 VGND X 0.03fF
C23 C X 0.00fF
C24 VPB a_29_53# 0.02fF
C25 VGND VPB 0.01fF
C26 X B 0.00fF
C27 VPWR X 0.07fF
C28 C VPB 0.01fF
C29 VPB B 0.03fF
C30 a_183_297# X 0.00fF
C31 VPWR VPB 0.05fF
C32 X a_111_297# 0.00fF
C33 a_29_53# A 0.26fF
C34 VGND A 0.01fF
C35 C A 0.03fF
C36 VGND a_29_53# 0.17fF
C37 B A 0.06fF
C38 C a_29_53# 0.06fF
C39 VPWR A 0.01fF
C40 VGND VNB 0.31fF
C41 X VNB 0.09fF
C42 A VNB 0.11fF
C43 C VNB 0.17fF
C44 B VNB 0.13fF
C45 VPWR VNB 0.28fF
C46 VPB VNB 0.52fF
C47 a_29_53# VNB 0.20fF
.ends

.subckt sky130_fd_sc_hd__inv_1 Y A VGND VPWR VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
C0 VGND A 0.03fF
C1 VGND VPB 0.01fF
C2 A VPB 0.02fF
C3 Y VPWR 0.11fF
C4 VGND Y 0.09fF
C5 A Y 0.02fF
C6 Y VPB 0.01fF
C7 VGND VPWR 0.04fF
C8 A VPWR 0.04fF
C9 VPB VPWR 0.04fF
C10 VGND VNB 0.25fF
C11 Y VNB 0.11fF
C12 VPWR VNB 0.24fF
C13 A VNB 0.19fF
C14 VPB VNB 0.34fF
.ends

.subckt sky130_fd_sc_hd__nor3_1 C Y A B VGND VPWR a_193_297# VNB VPB a_109_297#
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=3.445e+11p pd=3.66e+06u as=3.445e+11p ps=3.66e+06u w=650000u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 VGND VPB 0.01fF
C1 B Y 0.17fF
C2 B a_193_297# 0.00fF
C3 B VGND 0.01fF
C4 a_193_297# Y 0.01fF
C5 VPWR VPB 0.04fF
C6 VGND Y 0.12fF
C7 A VPB 0.02fF
C8 a_193_297# VGND 0.00fF
C9 B VPWR 0.01fF
C10 B A 0.06fF
C11 VPWR Y 0.13fF
C12 A Y 0.08fF
C13 a_193_297# VPWR 0.00fF
C14 a_193_297# A 0.00fF
C15 VGND VPWR 0.05fF
C16 VGND A 0.03fF
C17 C VPB 0.01fF
C18 A VPWR 0.03fF
C19 B C 0.08fF
C20 B a_109_297# 0.01fF
C21 C Y 0.07fF
C22 VGND C 0.01fF
C23 a_109_297# Y 0.00fF
C24 VGND a_109_297# 0.00fF
C25 C VPWR 0.01fF
C26 A C 0.00fF
C27 B VPB 0.01fF
C28 a_109_297# VPWR 0.00fF
C29 A a_109_297# 0.00fF
C30 VPB Y 0.01fF
C31 VGND VNB 0.27fF
C32 VPWR VNB 0.25fF
C33 Y VNB 0.10fF
C34 A VNB 0.19fF
C35 B VNB 0.08fF
C36 C VNB 0.15fF
C37 VPB VNB 0.43fF
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 Q RESET_B D CLK VGND VPWR a_1462_47# a_543_47# VNB
+ VPB a_651_413# a_193_47# a_805_47# a_448_47# a_639_47# a_1283_21# a_761_289# a_1108_47#
+ a_1217_47# a_1270_413# a_27_47#
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=1.0617e+12p pd=9.62e+06u as=0p ps=0u w=420000u l=150000u
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=1.2195e+12p ps=1.255e+07u w=1e+06u l=150000u
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X12 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_805_47# VPWR 0.00fF
C1 a_761_289# a_651_413# 0.09fF
C2 a_761_289# VGND 0.06fF
C3 a_1462_47# a_1283_21# 0.00fF
C4 a_639_47# VPWR 0.00fF
C5 Q a_27_47# 0.00fF
C6 a_448_47# a_27_47# 0.07fF
C7 a_761_289# a_1283_21# 0.00fF
C8 a_761_289# a_805_47# 0.00fF
C9 a_651_413# VGND 0.00fF
C10 VPWR Q 0.07fF
C11 a_448_47# VPWR 0.05fF
C12 a_761_289# a_639_47# 0.00fF
C13 a_651_413# a_1283_21# 0.00fF
C14 a_1462_47# Q 0.00fF
C15 a_1462_47# a_448_47# 0.00fF
C16 VGND a_1283_21# 0.18fF
C17 a_651_413# a_805_47# 0.00fF
C18 a_805_47# VGND 0.00fF
C19 a_1108_47# RESET_B 0.17fF
C20 a_761_289# Q 0.00fF
C21 a_761_289# a_448_47# 0.00fF
C22 a_651_413# a_639_47# 0.00fF
C23 a_639_47# VGND 0.00fF
C24 a_805_47# a_1283_21# 0.00fF
C25 a_543_47# RESET_B 0.15fF
C26 a_193_47# VPB 0.07fF
C27 a_639_47# a_1283_21# 0.00fF
C28 a_651_413# Q 0.00fF
C29 a_651_413# a_448_47# 0.00fF
C30 VGND Q 0.04fF
C31 a_448_47# VGND 0.06fF
C32 a_1108_47# a_27_47# 0.09fF
C33 Q a_1283_21# 0.04fF
C34 a_448_47# a_1283_21# 0.00fF
C35 a_193_47# a_1217_47# 0.00fF
C36 a_543_47# a_27_47# 0.05fF
C37 a_805_47# Q 0.00fF
C38 a_448_47# a_805_47# 0.00fF
C39 a_1108_47# VPWR 0.14fF
C40 VPB D 0.04fF
C41 VPB CLK 0.02fF
C42 a_639_47# Q 0.00fF
C43 a_639_47# a_448_47# 0.00fF
C44 a_1462_47# a_1108_47# 0.00fF
C45 a_543_47# VPWR 0.08fF
C46 a_193_47# D 0.15fF
C47 a_193_47# a_1270_413# 0.00fF
C48 a_193_47# CLK 0.00fF
C49 a_761_289# a_1108_47# 0.05fF
C50 a_1462_47# a_543_47# 0.00fF
C51 a_448_47# Q 0.00fF
C52 a_1217_47# D 0.00fF
C53 a_761_289# a_543_47# 0.15fF
C54 a_651_413# a_1108_47# 0.00fF
C55 a_1108_47# VGND 0.11fF
C56 a_1270_413# D 0.00fF
C57 CLK D 0.00fF
C58 a_651_413# a_543_47# 0.05fF
C59 a_1108_47# a_1283_21# 0.18fF
C60 a_543_47# VGND 0.10fF
C61 a_805_47# a_1108_47# 0.00fF
C62 a_543_47# a_1283_21# 0.00fF
C63 a_639_47# a_1108_47# 0.00fF
C64 a_543_47# a_805_47# 0.00fF
C65 a_639_47# a_543_47# 0.01fF
C66 a_1108_47# Q 0.00fF
C67 a_448_47# a_1108_47# 0.00fF
C68 VPB RESET_B 0.06fF
C69 a_543_47# Q 0.00fF
C70 a_448_47# a_543_47# 0.04fF
C71 a_193_47# RESET_B 0.02fF
C72 a_1217_47# RESET_B 0.00fF
C73 VPB a_27_47# 0.09fF
C74 a_193_47# a_27_47# 0.72fF
C75 D RESET_B 0.00fF
C76 a_1270_413# RESET_B 0.00fF
C77 VPB VPWR 0.19fF
C78 CLK RESET_B 0.00fF
C79 a_1217_47# a_27_47# 0.00fF
C80 a_193_47# VPWR 0.40fF
C81 a_543_47# a_1108_47# 0.00fF
C82 a_1462_47# a_193_47# 0.00fF
C83 a_1217_47# VPWR 0.00fF
C84 a_761_289# VPB 0.03fF
C85 D a_27_47# 0.09fF
C86 a_1270_413# a_27_47# 0.00fF
C87 CLK a_27_47# 0.19fF
C88 a_761_289# a_193_47# 0.12fF
C89 D VPWR 0.06fF
C90 a_651_413# VPB 0.01fF
C91 a_1270_413# VPWR 0.00fF
C92 a_761_289# a_1217_47# 0.00fF
C93 CLK VPWR 0.01fF
C94 VPB VGND 0.06fF
C95 a_1462_47# D 0.00fF
C96 a_651_413# a_193_47# 0.01fF
C97 a_193_47# VGND 0.05fF
C98 VPB a_1283_21# 0.05fF
C99 a_761_289# D 0.00fF
C100 a_1217_47# VGND 0.00fF
C101 a_761_289# a_1270_413# 0.00fF
C102 a_761_289# CLK 0.00fF
C103 a_193_47# a_1283_21# 0.04fF
C104 a_193_47# a_805_47# 0.00fF
C105 a_1217_47# a_1283_21# 0.00fF
C106 a_639_47# a_193_47# 0.00fF
C107 a_651_413# D 0.00fF
C108 D VGND 0.05fF
C109 a_651_413# a_1270_413# 0.00fF
C110 a_651_413# CLK 0.00fF
C111 VPB Q 0.01fF
C112 CLK VGND 0.01fF
C113 a_1270_413# VGND 0.00fF
C114 a_448_47# VPB 0.01fF
C115 D a_1283_21# 0.00fF
C116 a_193_47# Q 0.00fF
C117 a_448_47# a_193_47# 0.04fF
C118 a_1270_413# a_1283_21# 0.00fF
C119 CLK a_1283_21# 0.00fF
C120 a_805_47# D 0.00fF
C121 a_1217_47# Q 0.00fF
C122 a_448_47# a_1217_47# 0.00fF
C123 a_639_47# D 0.00fF
C124 RESET_B a_27_47# 0.33fF
C125 D Q 0.00fF
C126 a_448_47# D 0.12fF
C127 a_1270_413# Q 0.00fF
C128 a_448_47# CLK 0.00fF
C129 a_448_47# a_1270_413# 0.00fF
C130 RESET_B VPWR 0.06fF
C131 a_1462_47# RESET_B 0.00fF
C132 a_1108_47# VPB 0.04fF
C133 a_761_289# RESET_B 0.13fF
C134 a_193_47# a_1108_47# 0.10fF
C135 a_543_47# VPB 0.04fF
C136 VPWR a_27_47# 0.12fF
C137 a_1217_47# a_1108_47# 0.01fF
C138 a_543_47# a_193_47# 0.16fF
C139 a_1462_47# a_27_47# 0.00fF
C140 a_651_413# RESET_B 0.00fF
C141 RESET_B VGND 0.29fF
C142 a_543_47# a_1217_47# 0.00fF
C143 a_761_289# a_27_47# 0.04fF
C144 a_1108_47# D 0.00fF
C145 a_1462_47# VPWR 0.00fF
C146 a_1270_413# a_1108_47# 0.01fF
C147 RESET_B a_1283_21# 0.22fF
C148 a_1108_47# CLK 0.00fF
C149 a_805_47# RESET_B 0.00fF
C150 a_761_289# VPWR 0.08fF
C151 a_543_47# D 0.00fF
C152 a_543_47# a_1270_413# 0.00fF
C153 a_543_47# CLK 0.00fF
C154 a_651_413# a_27_47# 0.00fF
C155 a_639_47# RESET_B 0.00fF
C156 VGND a_27_47# 0.23fF
C157 a_761_289# a_1462_47# 0.00fF
C158 a_27_47# a_1283_21# 0.04fF
C159 a_651_413# VPWR 0.11fF
C160 RESET_B Q 0.00fF
C161 VPWR VGND 0.09fF
C162 a_448_47# RESET_B 0.00fF
C163 a_805_47# a_27_47# 0.00fF
C164 a_1462_47# VGND 0.00fF
C165 VPWR a_1283_21# 0.19fF
C166 a_639_47# a_27_47# 0.00fF
C167 Q VNB 0.09fF
C168 VGND VNB 1.04fF
C169 VPWR VNB 0.91fF
C170 RESET_B VNB 0.24fF
C171 D VNB 0.14fF
C172 CLK VNB 0.20fF
C173 VPB VNB 1.85fF
C174 a_651_413# VNB 0.00fF
C175 a_448_47# VNB 0.01fF
C176 a_1108_47# VNB 0.14fF
C177 a_1283_21# VNB 0.27fF
C178 a_543_47# VNB 0.14fF
C179 a_761_289# VNB 0.11fF
C180 a_193_47# VNB 0.25fF
C181 a_27_47# VNB 0.41fF
.ends

.subckt sky130_fd_sc_hd__a221oi_4 A2 Y C1 A1 B2 B1 VPWR VGND a_1241_47# VNB VPB a_453_47#
+ a_27_297# a_471_297#
X0 Y A1 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=1.053e+12p pd=1.104e+07u as=7.02e+11p ps=7.36e+06u w=650000u l=150000u
X1 a_453_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.027e+12p pd=8.36e+06u as=1.2935e+12p ps=1.308e+07u w=650000u l=150000u
X2 Y B1 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A1 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=1.89e+12p ps=1.778e+07u w=1e+06u l=150000u
X5 a_471_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.525e+12p pd=2.305e+07u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X6 Y B1 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND A2 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_453_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_471_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND B2 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_1241_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_27_297# B2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_453_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_1241_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_1241_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VPWR A2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_471_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_471_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_471_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR A1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_27_297# B1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND A2 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_471_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_27_297# B1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_1241_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 a_471_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 VPWR A1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_27_297# B2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_471_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_453_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 VGND B2 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 VGND VPWR 0.21fF
C1 VPWR C1 0.02fF
C2 Y VGND 0.45fF
C3 Y C1 0.19fF
C4 VGND VPB 0.05fF
C5 VGND B1 0.02fF
C6 VPB C1 0.05fF
C7 B1 C1 0.00fF
C8 A2 VPWR 0.04fF
C9 B2 a_1241_47# 0.00fF
C10 A2 Y 0.04fF
C11 A2 VPB 0.06fF
C12 A2 B1 0.00fF
C13 Y VPWR 0.02fF
C14 VPWR VPB 0.17fF
C15 B1 VPWR 0.02fF
C16 a_27_297# a_453_47# 0.00fF
C17 a_27_297# a_471_297# 0.38fF
C18 A1 a_27_297# 0.00fF
C19 Y VPB 0.02fF
C20 Y B1 0.18fF
C21 VGND B2 0.04fF
C22 B2 C1 0.04fF
C23 B1 VPB 0.05fF
C24 A2 B2 0.09fF
C25 a_471_297# a_453_47# 0.00fF
C26 A1 a_453_47# 0.00fF
C27 A1 a_471_297# 0.02fF
C28 VPWR B2 0.02fF
C29 Y B2 0.14fF
C30 B2 VPB 0.07fF
C31 B1 B2 0.32fF
C32 a_453_47# a_1241_47# 0.00fF
C33 a_471_297# a_1241_47# 0.00fF
C34 A1 a_1241_47# 0.02fF
C35 VGND a_27_297# 0.02fF
C36 a_27_297# C1 0.05fF
C37 A2 a_27_297# 0.00fF
C38 VGND a_453_47# 0.39fF
C39 a_453_47# C1 0.00fF
C40 VGND a_471_297# 0.02fF
C41 VGND A1 0.02fF
C42 a_471_297# C1 0.00fF
C43 A1 C1 0.00fF
C44 VPWR a_27_297# 0.19fF
C45 Y a_27_297# 0.44fF
C46 A2 a_453_47# 0.00fF
C47 A2 a_471_297# 0.45fF
C48 A2 A1 0.33fF
C49 a_27_297# VPB 0.02fF
C50 B1 a_27_297# 0.02fF
C51 VPWR a_453_47# 0.01fF
C52 VPWR a_471_297# 0.74fF
C53 A1 VPWR 0.04fF
C54 Y a_453_47# 0.23fF
C55 Y a_471_297# 0.01fF
C56 Y A1 0.10fF
C57 a_453_47# VPB 0.00fF
C58 B1 a_453_47# 0.02fF
C59 a_471_297# VPB 0.02fF
C60 B1 a_471_297# 0.02fF
C61 A1 VPB 0.05fF
C62 B1 A1 0.00fF
C63 VGND a_1241_47# 0.36fF
C64 a_1241_47# C1 0.00fF
C65 B2 a_27_297# 0.18fF
C66 A2 a_1241_47# 0.10fF
C67 B2 a_453_47# 0.01fF
C68 B2 a_471_297# 0.04fF
C69 A1 B2 0.00fF
C70 VPWR a_1241_47# 0.01fF
C71 VGND C1 0.06fF
C72 Y a_1241_47# 0.16fF
C73 a_1241_47# VPB 0.00fF
C74 B1 a_1241_47# 0.00fF
C75 A2 VGND 0.06fF
C76 A2 C1 0.00fF
C77 VGND VNB 1.09fF
C78 VPWR VNB 0.89fF
C79 Y VNB 0.06fF
C80 A1 VNB 0.32fF
C81 A2 VNB 0.39fF
C82 B1 VNB 0.32fF
C83 B2 VNB 0.39fF
C84 C1 VNB 0.39fF
C85 VPB VNB 1.93fF
C86 a_1241_47# VNB 0.01fF
C87 a_453_47# VNB 0.01fF
C88 a_471_297# VNB 0.06fF
C89 a_27_297# VNB 0.07fF
.ends

.subckt sky130_fd_sc_hd__nor2_1 B Y A VGND VPWR VNB VPB a_109_297#
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=3.38e+11p pd=3.64e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 Y A 0.03fF
C1 A VPWR 0.05fF
C2 B Y 0.06fF
C3 B VPWR 0.01fF
C4 B A 0.06fF
C5 Y a_109_297# 0.00fF
C6 a_109_297# VPWR 0.00fF
C7 Y VGND 0.14fF
C8 VGND VPWR 0.04fF
C9 VGND A 0.03fF
C10 B VGND 0.03fF
C11 VGND a_109_297# 0.00fF
C12 Y VPB 0.01fF
C13 VPB VPWR 0.04fF
C14 VPB A 0.02fF
C15 B VPB 0.02fF
C16 Y VPWR 0.08fF
C17 VGND VPB 0.01fF
C18 VGND VNB 0.27fF
C19 VPWR VNB 0.23fF
C20 Y VNB 0.08fF
C21 A VNB 0.16fF
C22 B VNB 0.15fF
C23 VPB VNB 0.34fF
.ends

.subckt sky130_fd_sc_hd__or2b_1 A B_N X VGND VPWR VNB VPB a_27_53# a_219_297# a_301_297#
X0 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=5.1875e+11p ps=4.32e+06u w=420000u l=150000u
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.057e+11p pd=4.04e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X3 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X4 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 VPB VGND 0.02fF
C1 A X 0.00fF
C2 X a_219_297# 0.06fF
C3 VPB X 0.01fF
C4 a_301_297# VPWR 0.00fF
C5 VGND X 0.03fF
C6 A B_N 0.00fF
C7 B_N a_219_297# 0.00fF
C8 VPB B_N 0.02fF
C9 A a_27_53# 0.11fF
C10 a_27_53# a_219_297# 0.08fF
C11 VPB a_27_53# 0.02fF
C12 VGND B_N 0.01fF
C13 VGND a_27_53# 0.10fF
C14 X B_N 0.00fF
C15 X a_27_53# 0.00fF
C16 A VPWR 0.14fF
C17 VPWR a_219_297# 0.06fF
C18 a_27_53# B_N 0.08fF
C19 A a_301_297# 0.00fF
C20 VPB VPWR 0.07fF
C21 a_301_297# a_219_297# 0.00fF
C22 VGND VPWR 0.07fF
C23 VGND a_301_297# 0.00fF
C24 X VPWR 0.07fF
C25 X a_301_297# 0.00fF
C26 B_N VPWR 0.03fF
C27 a_27_53# VPWR 0.03fF
C28 a_27_53# a_301_297# 0.00fF
C29 A a_219_297# 0.12fF
C30 VPB A 0.04fF
C31 VPB a_219_297# 0.02fF
C32 VGND A 0.01fF
C33 VGND a_219_297# 0.10fF
C34 VGND VNB 0.36fF
C35 X VNB 0.09fF
C36 B_N VNB 0.17fF
C37 A VNB 0.18fF
C38 VPWR VNB 0.36fF
C39 VPB VNB 0.60fF
C40 a_27_53# VNB 0.16fF
C41 a_219_297# VNB 0.15fF
.ends

.subckt sky130_fd_sc_hd__mux4_1 S0 A1 X S1 A2 A0 A3 VGND VPWR a_1290_413# a_757_363#
+ a_1478_413# a_277_47# VNB VPB a_750_97# a_27_413# a_923_363# a_193_47# a_834_97#
+ a_247_21# a_668_97# a_193_413# a_27_47#
X0 a_277_47# a_247_21# a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.226e+11p pd=2.74e+06u as=2.184e+11p ps=2.72e+06u w=420000u l=150000u
X1 VGND S0 a_247_21# VNB sky130_fd_pr__nfet_01v8 ad=6.142e+11p pd=7.3e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 a_834_97# a_247_21# a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=2.1715e+11p pd=2.72e+06u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X3 VGND A3 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.171e+11p ps=2.72e+06u w=420000u l=150000u
X4 a_1290_413# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=7.039e+11p ps=8e+06u w=420000u l=150000u
X5 a_834_97# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_750_97# S0 a_757_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.822e+11p pd=3.5e+06u as=2.171e+11p ps=2.72e+06u w=420000u l=150000u
X7 a_27_47# S0 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=2.184e+11p pd=2.72e+06u as=2.7965e+11p ps=3.21e+06u w=420000u l=150000u
X8 X a_1478_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9 VPWR A1 a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR S0 a_247_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.083e+11p ps=1.36e+06u w=420000u l=150000u
X11 X a_1478_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X12 a_193_47# A0 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13 a_750_97# a_1290_413# a_1478_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.84175e+11p ps=1.98e+06u w=420000u l=150000u
X14 a_1478_413# S1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_1290_413# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16 a_277_47# a_247_21# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_750_97# S0 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_923_363# a_247_21# a_750_97# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.8025e+11p pd=1.99e+06u as=0p ps=0u w=420000u l=150000u
X19 a_757_363# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR A3 a_923_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_277_47# a_1290_413# a_1478_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.0205e+11p ps=2.57e+06u w=420000u l=150000u
X22 a_193_413# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.171e+11p pd=2.72e+06u as=0p ps=0u w=420000u l=150000u
X23 a_193_413# S0 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_1478_413# S1 a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 A1 a_668_97# 0.00fF
C1 S1 X 0.00fF
C2 A3 A2 0.15fF
C3 a_27_413# A2 0.00fF
C4 A3 a_834_97# 0.04fF
C5 A2 a_1478_413# 0.00fF
C6 a_1478_413# a_834_97# 0.00fF
C7 a_277_47# A0 0.04fF
C8 VPB a_1290_413# 0.06fF
C9 a_247_21# a_668_97# 0.01fF
C10 A3 a_750_97# 0.02fF
C11 a_27_413# a_750_97# 0.00fF
C12 a_750_97# a_1478_413# 0.12fF
C13 S1 VPWR 0.03fF
C14 A2 A0 0.00fF
C15 a_757_363# A3 0.03fF
C16 a_757_363# a_27_413# 0.00fF
C17 A0 a_834_97# 0.00fF
C18 a_757_363# a_1478_413# 0.00fF
C19 A1 A3 0.00fF
C20 a_27_413# A1 0.03fF
C21 A1 a_1478_413# 0.00fF
C22 a_750_97# A0 0.00fF
C23 X VPB 0.01fF
C24 a_277_47# A2 0.00fF
C25 a_277_47# a_834_97# 0.02fF
C26 a_247_21# A3 0.06fF
C27 a_757_363# A0 0.00fF
C28 a_27_413# a_247_21# 0.00fF
C29 a_247_21# a_1478_413# 0.00fF
C30 A1 A0 0.14fF
C31 a_277_47# a_750_97# 0.23fF
C32 S1 VGND 0.03fF
C33 A2 a_834_97# 0.05fF
C34 VPB VPWR 0.20fF
C35 a_277_47# a_757_363# 0.00fF
C36 a_247_21# A0 0.06fF
C37 A2 a_750_97# 0.00fF
C38 S0 a_193_413# 0.01fF
C39 a_277_47# A1 0.00fF
C40 a_750_97# a_834_97# 0.03fF
C41 a_193_47# a_1290_413# 0.00fF
C42 a_757_363# A2 0.04fF
C43 a_757_363# a_834_97# 0.01fF
C44 a_277_47# a_247_21# 0.31fF
C45 A1 A2 0.00fF
C46 a_27_47# S0 0.00fF
C47 A1 a_834_97# 0.00fF
C48 a_757_363# a_750_97# 0.10fF
C49 X a_1290_413# 0.00fF
C50 VGND VPB 0.06fF
C51 A1 a_750_97# 0.00fF
C52 a_247_21# A2 0.00fF
C53 a_247_21# a_834_97# 0.02fF
C54 a_757_363# A1 0.00fF
C55 a_27_47# a_668_97# 0.00fF
C56 a_247_21# a_750_97# 0.09fF
C57 a_1290_413# VPWR 0.08fF
C58 a_923_363# a_1290_413# 0.00fF
C59 a_757_363# a_247_21# 0.01fF
C60 A3 a_193_413# 0.00fF
C61 a_27_413# a_193_413# 0.07fF
C62 a_193_413# a_1478_413# 0.00fF
C63 a_247_21# A1 0.00fF
C64 a_193_47# VPWR 0.00fF
C65 a_27_47# A3 0.00fF
C66 a_27_413# a_27_47# 0.01fF
C67 a_27_47# a_1478_413# 0.00fF
C68 a_193_413# A0 0.00fF
C69 X VPWR 0.04fF
C70 VGND a_1290_413# 0.07fF
C71 X a_923_363# 0.00fF
C72 S1 S0 0.00fF
C73 VGND a_193_47# 0.00fF
C74 a_27_47# A0 0.03fF
C75 a_277_47# a_193_413# 0.06fF
C76 a_923_363# VPWR 0.00fF
C77 A2 a_193_413# 0.00fF
C78 X VGND 0.04fF
C79 a_277_47# a_27_47# 0.07fF
C80 S1 a_668_97# 0.00fF
C81 a_750_97# a_193_413# 0.00fF
C82 a_27_47# A2 0.00fF
C83 S0 VPB 0.11fF
C84 a_27_47# a_834_97# 0.00fF
C85 VGND VPWR 0.09fF
C86 a_757_363# a_193_413# 0.00fF
C87 VGND a_923_363# 0.00fF
C88 A1 a_193_413# 0.00fF
C89 a_27_47# a_750_97# 0.00fF
C90 S1 A3 0.00fF
C91 a_27_413# S1 0.00fF
C92 S1 a_1478_413# 0.00fF
C93 VPB a_668_97# 0.00fF
C94 a_247_21# a_193_413# 0.07fF
C95 a_27_47# A1 0.03fF
C96 S1 A0 0.00fF
C97 a_247_21# a_27_47# 0.03fF
C98 S0 a_1290_413# 0.00fF
C99 A3 VPB 0.03fF
C100 a_27_413# VPB 0.01fF
C101 a_277_47# S1 0.01fF
C102 VPB a_1478_413# 0.04fF
C103 S1 A2 0.05fF
C104 S1 a_834_97# 0.00fF
C105 VPB A0 0.03fF
C106 a_1290_413# a_668_97# 0.00fF
C107 S1 a_750_97# 0.01fF
C108 X S0 0.00fF
C109 a_193_47# a_668_97# 0.00fF
C110 a_757_363# S1 0.00fF
C111 a_277_47# VPB 0.02fF
C112 S1 A1 0.00fF
C113 S0 VPWR 0.05fF
C114 X a_668_97# 0.00fF
C115 A3 a_1290_413# 0.00fF
C116 a_923_363# S0 0.00fF
C117 a_27_413# a_1290_413# 0.00fF
C118 A2 VPB 0.02fF
C119 a_1290_413# a_1478_413# 0.07fF
C120 VPB a_834_97# 0.01fF
C121 a_247_21# S1 0.00fF
C122 a_27_47# a_193_413# 0.00fF
C123 VPB a_750_97# 0.04fF
C124 a_27_413# a_193_47# 0.00fF
C125 a_193_47# a_1478_413# 0.00fF
C126 a_1290_413# A0 0.00fF
C127 VPWR a_668_97# 0.00fF
C128 a_757_363# VPB 0.02fF
C129 a_923_363# a_668_97# 0.00fF
C130 A1 VPB 0.02fF
C131 X A3 0.00fF
C132 VGND S0 0.03fF
C133 a_27_413# X 0.00fF
C134 X a_1478_413# 0.07fF
C135 a_193_47# A0 0.00fF
C136 a_277_47# a_1290_413# 0.35fF
C137 a_247_21# VPB 0.07fF
C138 A3 VPWR 0.01fF
C139 a_27_413# VPWR 0.07fF
C140 a_277_47# a_193_47# 0.00fF
C141 VGND a_668_97# 0.18fF
C142 VPWR a_1478_413# 0.16fF
C143 A2 a_1290_413# 0.00fF
C144 a_923_363# A3 0.00fF
C145 a_27_413# a_923_363# 0.00fF
C146 a_1290_413# a_834_97# 0.01fF
C147 a_923_363# a_1478_413# 0.00fF
C148 a_750_97# a_1290_413# 0.13fF
C149 a_193_47# a_834_97# 0.00fF
C150 a_277_47# X 0.00fF
C151 VPWR A0 0.01fF
C152 a_757_363# a_1290_413# 0.01fF
C153 a_193_47# a_750_97# 0.00fF
C154 A1 a_1290_413# 0.00fF
C155 S1 a_193_413# 0.00fF
C156 X A2 0.00fF
C157 VGND A3 0.01fF
C158 a_27_413# VGND 0.00fF
C159 X a_834_97# 0.00fF
C160 VGND a_1478_413# 0.15fF
C161 a_277_47# VPWR 0.05fF
C162 a_277_47# a_923_363# 0.00fF
C163 X a_750_97# 0.00fF
C164 a_247_21# a_1290_413# 0.01fF
C165 S1 a_27_47# 0.00fF
C166 VGND A0 0.01fF
C167 a_757_363# X 0.00fF
C168 A2 VPWR 0.01fF
C169 VPWR a_834_97# 0.00fF
C170 a_247_21# a_193_47# 0.00fF
C171 a_923_363# a_834_97# 0.00fF
C172 a_750_97# VPWR 0.23fF
C173 a_923_363# a_750_97# 0.00fF
C174 VPB a_193_413# 0.01fF
C175 a_277_47# VGND 0.42fF
C176 a_247_21# X 0.00fF
C177 a_757_363# VPWR 0.20fF
C178 a_757_363# a_923_363# 0.01fF
C179 A1 VPWR 0.01fF
C180 a_27_47# VPB 0.01fF
C181 VGND A2 0.01fF
C182 VGND a_834_97# 0.08fF
C183 a_247_21# VPWR 0.13fF
C184 VGND a_750_97# 0.05fF
C185 a_247_21# a_923_363# 0.00fF
C186 S0 a_668_97# 0.02fF
C187 a_757_363# VGND 0.00fF
C188 VGND A1 0.01fF
C189 a_193_413# a_1290_413# 0.00fF
C190 a_247_21# VGND 0.08fF
C191 S0 A3 0.00fF
C192 a_27_413# S0 0.00fF
C193 a_193_47# a_193_413# 0.00fF
C194 S0 a_1478_413# 0.00fF
C195 a_27_47# a_1290_413# 0.00fF
C196 a_27_47# a_193_47# 0.00fF
C197 X a_193_413# 0.00fF
C198 S0 A0 0.00fF
C199 A3 a_668_97# 0.00fF
C200 S1 VPB 0.06fF
C201 a_668_97# a_1478_413# 0.00fF
C202 X a_27_47# 0.00fF
C203 a_277_47# S0 0.01fF
C204 a_193_413# VPWR 0.15fF
C205 A0 a_668_97# 0.00fF
C206 a_923_363# a_193_413# 0.00fF
C207 S0 A2 0.00fF
C208 a_27_413# A3 0.00fF
C209 S0 a_834_97# 0.00fF
C210 A3 a_1478_413# 0.00fF
C211 a_27_413# a_1478_413# 0.00fF
C212 a_27_47# VPWR 0.01fF
C213 a_277_47# a_668_97# 0.00fF
C214 S0 a_750_97# 0.05fF
C215 VGND a_193_413# 0.00fF
C216 A3 A0 0.00fF
C217 a_27_413# A0 0.06fF
C218 a_757_363# S0 0.02fF
C219 A0 a_1478_413# 0.00fF
C220 S1 a_1290_413# 0.12fF
C221 A2 a_668_97# 0.00fF
C222 a_668_97# a_834_97# 0.06fF
C223 A1 S0 0.00fF
C224 a_750_97# a_668_97# 0.06fF
C225 VGND a_27_47# 0.18fF
C226 a_277_47# A3 0.00fF
C227 a_277_47# a_27_413# 0.05fF
C228 a_277_47# a_1478_413# 0.08fF
C229 a_247_21# S0 0.28fF
C230 a_757_363# a_668_97# 0.00fF
C231 VGND VNB 1.09fF
C232 X VNB 0.09fF
C233 S1 VNB 0.30fF
C234 A2 VNB 0.08fF
C235 A3 VNB 0.10fF
C236 S0 VNB 0.42fF
C237 VPWR VNB 0.95fF
C238 A0 VNB 0.08fF
C239 A1 VNB 0.19fF
C240 VPB VNB 1.93fF
C241 a_834_97# VNB 0.03fF
C242 a_668_97# VNB 0.01fF
C243 a_27_47# VNB 0.05fF
C244 a_1478_413# VNB 0.16fF
C245 a_1290_413# VNB 0.23fF
C246 a_750_97# VNB 0.06fF
C247 a_757_363# VNB 0.01fF
C248 a_277_47# VNB 0.09fF
C249 a_247_21# VNB 0.28fF
C250 a_193_413# VNB 0.01fF
C251 a_27_413# VNB 0.04fF
.ends

.subckt sky130_fd_sc_hd__nor3_2 C Y A B VGND VPWR VNB VPB a_281_297# a_27_297#
X0 Y C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=7.9e+11p ps=7.58e+06u w=1e+06u l=150000u
X1 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.3e+11p ps=7.66e+06u w=1e+06u l=150000u
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=8.6125e+11p ps=9.15e+06u w=650000u l=150000u
X3 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_281_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 VPB A 0.02fF
C1 VPB a_27_297# 0.01fF
C2 VPB B 0.02fF
C3 Y a_281_297# 0.12fF
C4 A VGND 0.03fF
C5 VGND a_27_297# 0.01fF
C6 Y VPWR 0.01fF
C7 A a_27_297# 0.07fF
C8 VPB a_281_297# 0.01fF
C9 Y C 0.12fF
C10 B VGND 0.01fF
C11 A B 0.07fF
C12 B a_27_297# 0.09fF
C13 VPB VPWR 0.07fF
C14 VPB C 0.03fF
C15 VGND a_281_297# 0.01fF
C16 A a_281_297# 0.00fF
C17 a_281_297# a_27_297# 0.17fF
C18 VGND VPWR 0.08fF
C19 B a_281_297# 0.01fF
C20 A VPWR 0.01fF
C21 VGND C 0.01fF
C22 A C 0.00fF
C23 a_27_297# VPWR 0.21fF
C24 a_27_297# C 0.01fF
C25 B VPWR 0.01fF
C26 VPB Y 0.01fF
C27 B C 0.03fF
C28 a_281_297# VPWR 0.18fF
C29 Y VGND 0.46fF
C30 a_281_297# C 0.04fF
C31 A Y 0.05fF
C32 Y a_27_297# 0.01fF
C33 C VPWR 0.01fF
C34 B Y 0.12fF
C35 VPB VGND 0.02fF
C36 VGND VNB 0.49fF
C37 Y VNB 0.09fF
C38 VPWR VNB 0.38fF
C39 C VNB 0.20fF
C40 B VNB 0.16fF
C41 A VNB 0.21fF
C42 VPB VNB 0.78fF
C43 a_281_297# VNB 0.04fF
C44 a_27_297# VNB 0.05fF
.ends

.subckt sky130_fd_sc_hd__nand3b_1 B C A_N Y VGND VPWR VNB VPB a_53_93# a_232_47# a_316_47#
X0 Y a_53_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=5.5e+11p pd=5.1e+06u as=6.765e+11p ps=5.44e+06u w=1e+06u l=150000u
X1 a_232_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=2.005e+11p ps=1.97e+06u w=650000u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A_N a_53_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X4 VGND A_N a_53_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X5 a_316_47# B a_232_47# VNB sky130_fd_pr__nfet_01v8 ad=2.5025e+11p pd=2.07e+06u as=0p ps=0u w=650000u l=150000u
X6 Y a_53_93# a_316_47# VNB sky130_fd_pr__nfet_01v8 ad=1.82e+11p pd=1.86e+06u as=0p ps=0u w=650000u l=150000u
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 VPB VGND 0.02fF
C1 C B 0.08fF
C2 VPWR Y 0.30fF
C3 Y a_53_93# 0.09fF
C4 VPB Y 0.02fF
C5 a_316_47# B 0.00fF
C6 VGND Y 0.06fF
C7 VPWR A_N 0.01fF
C8 A_N a_53_93# 0.08fF
C9 VPB A_N 0.02fF
C10 VPWR a_232_47# 0.00fF
C11 a_232_47# a_53_93# 0.00fF
C12 VGND A_N 0.00fF
C13 VGND a_232_47# 0.00fF
C14 Y A_N 0.00fF
C15 Y a_232_47# 0.00fF
C16 VPWR C 0.01fF
C17 C a_53_93# 0.04fF
C18 VPB C 0.01fF
C19 VGND C 0.01fF
C20 VPWR B 0.01fF
C21 B a_53_93# 0.11fF
C22 VPWR a_316_47# 0.00fF
C23 VPB B 0.01fF
C24 a_316_47# a_53_93# 0.00fF
C25 VGND B 0.01fF
C26 Y C 0.01fF
C27 VGND a_316_47# 0.00fF
C28 Y B 0.05fF
C29 Y a_316_47# 0.00fF
C30 C A_N 0.06fF
C31 a_232_47# C 0.00fF
C32 A_N B 0.00fF
C33 a_232_47# B 0.00fF
C34 VPWR a_53_93# 0.05fF
C35 VPB VPWR 0.06fF
C36 VPB a_53_93# 0.02fF
C37 VGND VPWR 0.06fF
C38 VGND a_53_93# 0.12fF
C39 VGND VNB 0.36fF
C40 Y VNB 0.12fF
C41 A_N VNB 0.14fF
C42 VPWR VNB 0.33fF
C43 B VNB 0.08fF
C44 C VNB 0.09fF
C45 VPB VNB 0.60fF
C46 a_53_93# VNB 0.21fF
.ends

.subckt sky130_fd_sc_hd__or3b_2 A B C_N X VPWR VGND VNB VPB a_472_297# a_388_297#
+ a_176_21# a_27_47#
X0 a_388_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=5.88e+11p ps=5.35e+06u w=420000u l=150000u
X1 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=5.1765e+11p pd=5.33e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X5 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_176_21# a_27_47# a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X8 a_472_297# B a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
C0 a_176_21# VGND 0.17fF
C1 C_N VGND 0.01fF
C2 a_388_297# A 0.00fF
C3 a_176_21# VPB 0.03fF
C4 VPB C_N 0.03fF
C5 a_472_297# VGND 0.00fF
C6 a_176_21# a_388_297# 0.00fF
C7 a_388_297# C_N 0.00fF
C8 VPB VGND 0.02fF
C9 B VPWR 0.09fF
C10 a_27_47# A 0.11fF
C11 a_388_297# VGND 0.00fF
C12 X A 0.01fF
C13 a_176_21# a_27_47# 0.12fF
C14 a_27_47# C_N 0.10fF
C15 a_176_21# X 0.08fF
C16 X C_N 0.00fF
C17 a_472_297# a_27_47# 0.00fF
C18 a_472_297# X 0.00fF
C19 a_27_47# VGND 0.07fF
C20 VPB a_27_47# 0.03fF
C21 X VGND 0.07fF
C22 X VPB 0.00fF
C23 a_388_297# a_27_47# 0.00fF
C24 a_388_297# X 0.00fF
C25 VPWR A 0.01fF
C26 B A 0.06fF
C27 a_176_21# VPWR 0.02fF
C28 VPWR C_N 0.01fF
C29 X a_27_47# 0.11fF
C30 a_176_21# B 0.03fF
C31 B C_N 0.00fF
C32 a_472_297# VPWR 0.00fF
C33 a_472_297# B 0.00fF
C34 VPWR VGND 0.07fF
C35 VPB VPWR 0.07fF
C36 B VGND 0.01fF
C37 B VPB 0.03fF
C38 a_388_297# VPWR 0.00fF
C39 a_388_297# B 0.00fF
C40 a_27_47# VPWR 0.12fF
C41 B a_27_47# 0.14fF
C42 X VPWR 0.00fF
C43 X B 0.00fF
C44 a_176_21# A 0.10fF
C45 A C_N 0.00fF
C46 a_176_21# C_N 0.04fF
C47 a_472_297# A 0.00fF
C48 A VGND 0.01fF
C49 VPB A 0.02fF
C50 a_472_297# a_176_21# 0.00fF
C51 a_472_297# C_N 0.00fF
C52 VGND VNB 0.40fF
C53 A VNB 0.10fF
C54 B VNB 0.13fF
C55 X VNB 0.01fF
C56 C_N VNB 0.22fF
C57 VPWR VNB 0.36fF
C58 VPB VNB 0.69fF
C59 a_27_47# VNB 0.22fF
C60 a_176_21# VNB 0.26fF
.ends

.subckt sky130_fd_sc_hd__o2111a_2 D1 C1 A2 A1 B1 X VGND VPWR VNB a_386_47# VPB a_80_21#
+ a_674_297# a_566_47# a_458_47#
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=1.65e+12p pd=1.13e+07u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X1 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_80_21# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=6.7e+11p pd=5.34e+06u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=5.98e+11p pd=5.74e+06u as=1.82e+11p ps=1.86e+06u w=650000u l=150000u
X4 VPWR C1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_674_297# A2 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X8 a_386_47# D1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=1.7225e+11p ps=1.83e+06u w=650000u l=150000u
X9 VPWR A1 a_674_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_566_47# B1 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=4.2575e+11p pd=3.91e+06u as=2.535e+11p ps=2.08e+06u w=650000u l=150000u
X11 VGND A2 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_566_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_458_47# C1 a_386_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 D1 a_566_47# 0.00fF
C1 a_80_21# a_566_47# 0.00fF
C2 D1 X 0.00fF
C3 X a_80_21# 0.13fF
C4 VPWR D1 0.01fF
C5 VGND A1 0.02fF
C6 VPWR a_80_21# 0.27fF
C7 A2 a_566_47# 0.05fF
C8 D1 B1 0.00fF
C9 B1 a_80_21# 0.06fF
C10 A2 X 0.00fF
C11 A2 VPWR 0.09fF
C12 X a_566_47# 0.00fF
C13 VPWR a_566_47# 0.01fF
C14 A2 B1 0.08fF
C15 VPWR X 0.13fF
C16 C1 a_458_47# 0.00fF
C17 B1 a_566_47# 0.02fF
C18 B1 X 0.00fF
C19 A1 VPB 0.03fF
C20 VPWR B1 0.01fF
C21 D1 C1 0.10fF
C22 C1 a_80_21# 0.09fF
C23 D1 a_674_297# 0.00fF
C24 a_674_297# a_80_21# 0.00fF
C25 A2 C1 0.00fF
C26 A2 a_674_297# 0.01fF
C27 C1 a_566_47# 0.02fF
C28 VGND a_458_47# 0.00fF
C29 X C1 0.00fF
C30 a_674_297# a_566_47# 0.00fF
C31 VPWR C1 0.01fF
C32 a_674_297# X 0.00fF
C33 D1 VGND 0.01fF
C34 VGND a_80_21# 0.12fF
C35 VPWR a_674_297# 0.00fF
C36 B1 C1 0.08fF
C37 B1 a_674_297# 0.00fF
C38 A2 VGND 0.01fF
C39 VGND a_566_47# 0.13fF
C40 VGND X 0.10fF
C41 VPWR VGND 0.12fF
C42 D1 VPB 0.01fF
C43 VPB a_80_21# 0.04fF
C44 B1 VGND 0.01fF
C45 a_674_297# C1 0.00fF
C46 a_386_47# a_80_21# 0.00fF
C47 A2 VPB 0.02fF
C48 D1 A1 0.00fF
C49 VPB a_566_47# 0.00fF
C50 A1 a_80_21# 0.00fF
C51 X VPB 0.00fF
C52 a_386_47# a_566_47# 0.00fF
C53 VPWR VPB 0.10fF
C54 a_386_47# X 0.00fF
C55 VGND C1 0.04fF
C56 VPWR a_386_47# 0.00fF
C57 A2 A1 0.07fF
C58 B1 VPB 0.01fF
C59 VGND a_674_297# 0.00fF
C60 A1 a_566_47# 0.04fF
C61 A1 X 0.00fF
C62 VPWR A1 0.10fF
C63 B1 A1 0.00fF
C64 C1 VPB 0.01fF
C65 a_386_47# C1 0.00fF
C66 a_458_47# a_80_21# 0.00fF
C67 A1 C1 0.00fF
C68 D1 a_80_21# 0.15fF
C69 a_674_297# A1 0.00fF
C70 VGND VPB 0.03fF
C71 a_458_47# a_566_47# 0.00fF
C72 X a_458_47# 0.00fF
C73 VGND a_386_47# 0.00fF
C74 A2 D1 0.00fF
C75 A2 a_80_21# 0.03fF
C76 VPWR a_458_47# 0.00fF
C77 VGND VNB 0.57fF
C78 X VNB 0.03fF
C79 VPWR VNB 0.52fF
C80 A1 VNB 0.20fF
C81 A2 VNB 0.08fF
C82 B1 VNB 0.08fF
C83 C1 VNB 0.09fF
C84 D1 VNB 0.09fF
C85 VPB VNB 0.96fF
C86 a_566_47# VNB 0.04fF
C87 a_80_21# VNB 0.25fF
.ends

.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N Q RESET_B D VGND VPWR a_1462_47# a_543_47#
+ VNB VPB a_651_413# a_193_47# a_805_47# a_448_47# a_639_47# a_1283_21# a_761_289#
+ a_1108_47# a_1217_47# a_1270_413# a_27_47#
X0 a_1217_47# a_193_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X2 a_1108_47# a_27_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X4 a_651_413# a_193_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=1.0617e+12p pd=9.62e+06u as=0p ps=0u w=420000u l=150000u
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=1.2195e+12p ps=1.255e+07u w=1e+06u l=150000u
X7 VPWR CLK_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X11 a_1108_47# a_193_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X12 a_543_47# a_193_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_27_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X18 a_1270_413# a_27_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X23 a_639_47# a_27_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND CLK_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_1283_21# D 0.00fF
C1 a_1462_47# a_761_289# 0.00fF
C2 RESET_B a_805_47# 0.00fF
C3 a_193_47# a_805_47# 0.00fF
C4 Q a_27_47# 0.00fF
C5 a_651_413# a_1108_47# 0.00fF
C6 a_1108_47# VPB 0.04fF
C7 D RESET_B 0.00fF
C8 a_193_47# D 0.17fF
C9 a_1283_21# a_651_413# 0.00fF
C10 a_448_47# a_543_47# 0.04fF
C11 a_1283_21# VPB 0.05fF
C12 a_1462_47# a_1108_47# 0.00fF
C13 Q a_1270_413# 0.00fF
C14 a_1462_47# a_1283_21# 0.00fF
C15 a_761_289# a_1217_47# 0.00fF
C16 a_651_413# RESET_B 0.00fF
C17 a_651_413# a_193_47# 0.00fF
C18 RESET_B VPB 0.06fF
C19 a_193_47# VPB 0.06fF
C20 a_761_289# a_1108_47# 0.05fF
C21 a_1462_47# RESET_B 0.00fF
C22 a_1462_47# a_193_47# 0.00fF
C23 a_761_289# a_1283_21# 0.00fF
C24 VPWR a_805_47# 0.00fF
C25 a_1108_47# a_1217_47# 0.01fF
C26 D VPWR 0.06fF
C27 a_1283_21# a_1217_47# 0.00fF
C28 a_761_289# RESET_B 0.13fF
C29 a_761_289# a_193_47# 0.04fF
C30 VGND a_639_47# 0.00fF
C31 a_1283_21# a_1108_47# 0.18fF
C32 a_27_47# a_805_47# 0.00fF
C33 D a_27_47# 0.07fF
C34 a_651_413# VPWR 0.11fF
C35 RESET_B a_1217_47# 0.00fF
C36 VPWR VPB 0.19fF
C37 a_193_47# a_1217_47# 0.00fF
C38 a_448_47# Q 0.00fF
C39 RESET_B a_1108_47# 0.17fF
C40 a_193_47# a_1108_47# 0.09fF
C41 CLK_N D 0.00fF
C42 a_1462_47# VPWR 0.00fF
C43 a_1270_413# D 0.00fF
C44 a_1283_21# RESET_B 0.22fF
C45 a_1283_21# a_193_47# 0.04fF
C46 a_651_413# a_27_47# 0.01fF
C47 a_27_47# VPB 0.09fF
C48 VGND a_543_47# 0.10fF
C49 a_639_47# a_543_47# 0.01fF
C50 a_651_413# CLK_N 0.00fF
C51 a_1462_47# a_27_47# 0.00fF
C52 a_761_289# VPWR 0.08fF
C53 CLK_N VPB 0.02fF
C54 a_193_47# RESET_B 0.33fF
C55 a_651_413# a_1270_413# 0.00fF
C56 VPWR a_1217_47# 0.00fF
C57 a_761_289# a_27_47# 0.12fF
C58 VPWR a_1108_47# 0.14fF
C59 a_1283_21# VPWR 0.19fF
C60 a_761_289# CLK_N 0.00fF
C61 a_761_289# a_1270_413# 0.00fF
C62 a_27_47# a_1217_47# 0.00fF
C63 a_448_47# a_805_47# 0.00fF
C64 a_448_47# D 0.12fF
C65 a_1108_47# a_27_47# 0.10fF
C66 RESET_B VPWR 0.06fF
C67 a_193_47# VPWR 0.06fF
C68 a_1283_21# a_27_47# 0.04fF
C69 CLK_N a_1108_47# 0.00fF
C70 VGND Q 0.04fF
C71 a_1270_413# a_1108_47# 0.01fF
C72 Q a_639_47# 0.00fF
C73 a_1283_21# CLK_N 0.00fF
C74 a_651_413# a_448_47# 0.00fF
C75 a_448_47# VPB 0.01fF
C76 a_1283_21# a_1270_413# 0.00fF
C77 RESET_B a_27_47# 0.02fF
C78 a_193_47# a_27_47# 0.72fF
C79 a_1462_47# a_448_47# 0.00fF
C80 CLK_N RESET_B 0.00fF
C81 a_193_47# CLK_N 0.00fF
C82 a_1270_413# RESET_B 0.00fF
C83 a_193_47# a_1270_413# 0.00fF
C84 Q a_543_47# 0.00fF
C85 a_761_289# a_448_47# 0.00fF
C86 a_448_47# a_1217_47# 0.00fF
C87 VPWR a_27_47# 0.46fF
C88 a_448_47# a_1108_47# 0.00fF
C89 VGND a_805_47# 0.00fF
C90 CLK_N VPWR 0.01fF
C91 VGND D 0.05fF
C92 a_1283_21# a_448_47# 0.00fF
C93 a_639_47# D 0.00fF
C94 a_1270_413# VPWR 0.00fF
C95 a_448_47# RESET_B 0.00fF
C96 a_193_47# a_448_47# 0.08fF
C97 CLK_N a_27_47# 0.18fF
C98 a_651_413# VGND 0.00fF
C99 a_1270_413# a_27_47# 0.00fF
C100 VGND VPB 0.06fF
C101 a_651_413# a_639_47# 0.00fF
C102 a_543_47# a_805_47# 0.00fF
C103 a_1462_47# VGND 0.00fF
C104 a_543_47# D 0.00fF
C105 a_761_289# VGND 0.06fF
C106 a_761_289# a_639_47# 0.00fF
C107 a_651_413# a_543_47# 0.05fF
C108 a_543_47# VPB 0.04fF
C109 a_448_47# VPWR 0.05fF
C110 VGND a_1217_47# 0.00fF
C111 a_1462_47# a_543_47# 0.00fF
C112 VGND a_1108_47# 0.11fF
C113 a_639_47# a_1108_47# 0.00fF
C114 a_448_47# a_27_47# 0.04fF
C115 a_1283_21# VGND 0.18fF
C116 a_1283_21# a_639_47# 0.00fF
C117 a_761_289# a_543_47# 0.15fF
C118 a_448_47# CLK_N 0.00fF
C119 Q a_805_47# 0.00fF
C120 a_448_47# a_1270_413# 0.00fF
C121 Q D 0.00fF
C122 VGND RESET_B 0.29fF
C123 a_193_47# VGND 0.17fF
C124 a_639_47# RESET_B 0.00fF
C125 a_193_47# a_639_47# 0.00fF
C126 a_543_47# a_1217_47# 0.00fF
C127 a_543_47# a_1108_47# 0.00fF
C128 a_1283_21# a_543_47# 0.00fF
C129 a_651_413# Q 0.00fF
C130 Q VPB 0.01fF
C131 a_1462_47# Q 0.00fF
C132 a_543_47# RESET_B 0.15fF
C133 a_193_47# a_543_47# 0.05fF
C134 VGND VPWR 0.09fF
C135 a_639_47# VPWR 0.00fF
C136 a_761_289# Q 0.00fF
C137 D a_805_47# 0.00fF
C138 VGND a_27_47# 0.11fF
C139 Q a_1217_47# 0.00fF
C140 a_639_47# a_27_47# 0.00fF
C141 Q a_1108_47# 0.00fF
C142 CLK_N VGND 0.01fF
C143 VGND a_1270_413# 0.00fF
C144 a_543_47# VPWR 0.08fF
C145 a_1283_21# Q 0.04fF
C146 a_651_413# a_805_47# 0.00fF
C147 a_651_413# D 0.00fF
C148 D VPB 0.04fF
C149 Q RESET_B 0.00fF
C150 a_193_47# Q 0.00fF
C151 a_1462_47# D 0.00fF
C152 a_543_47# a_27_47# 0.16fF
C153 CLK_N a_543_47# 0.00fF
C154 a_651_413# VPB 0.01fF
C155 a_1270_413# a_543_47# 0.00fF
C156 a_761_289# a_805_47# 0.00fF
C157 a_761_289# D 0.00fF
C158 D a_1217_47# 0.00fF
C159 a_448_47# VGND 0.06fF
C160 a_1108_47# a_805_47# 0.00fF
C161 a_448_47# a_639_47# 0.00fF
C162 a_761_289# a_651_413# 0.09fF
C163 D a_1108_47# 0.00fF
C164 Q VPWR 0.07fF
C165 a_761_289# VPB 0.03fF
C166 a_1283_21# a_805_47# 0.00fF
C167 Q VNB 0.09fF
C168 VGND VNB 1.04fF
C169 VPWR VNB 0.91fF
C170 RESET_B VNB 0.24fF
C171 D VNB 0.14fF
C172 CLK_N VNB 0.20fF
C173 VPB VNB 1.85fF
C174 a_651_413# VNB 0.00fF
C175 a_448_47# VNB 0.01fF
C176 a_1108_47# VNB 0.14fF
C177 a_1283_21# VNB 0.27fF
C178 a_543_47# VNB 0.14fF
C179 a_761_289# VNB 0.11fF
C180 a_193_47# VNB 0.25fF
C181 a_27_47# VNB 0.41fF
.ends

.subckt SLC VOUT INB IN a_919_243# a_1235_416# a_264_22# VGND a_438_293# VNB VPB vpwr
X0 VGND IN a_264_22# VNB sky130_fd_pr__nfet_01v8_lvt ad=1.8755e+12p pd=2.064e+07u as=7.25e+11p ps=7.9e+06u w=500000u l=150000u
X1 a_264_22# IN VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2 a_919_243# INB VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=7.25e+11p pd=7.9e+06u as=0p ps=0u w=500000u l=150000u
X3 a_264_22# IN VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4 VGND INB a_919_243# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5 VGND INB a_919_243# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6 a_438_293# a_264_22# a_264_22# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.044e+11p pd=1.3e+06u as=9.72e+10p ps=1.26e+06u w=360000u l=150000u
X7 a_264_22# IN VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X8 a_264_22# IN VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X9 vpwr a_438_293# VOUT VPB sky130_fd_pr__pfet_01v8_hvt ad=4.819e+11p pd=5.67e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=150000u
X10 VGND a_264_22# VOUT VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X11 VGND IN a_264_22# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X12 VGND INB a_919_243# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X13 VGND IN a_264_22# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X14 a_919_243# INB VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X15 a_919_243# INB VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X16 a_1235_416# a_264_22# vpwr VPB sky130_fd_pr__pfet_01v8_hvt ad=1.044e+11p pd=1.3e+06u as=0p ps=0u w=360000u l=150000u
X17 VGND INB a_919_243# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X18 VGND IN a_264_22# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X19 VGND IN a_264_22# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X20 a_919_243# INB VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X21 VOUT a_438_293# vpwr VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X22 vpwr a_919_243# a_438_293# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23 a_264_22# IN VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X24 a_919_243# INB VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X25 VGND INB a_919_243# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X26 a_919_243# a_919_243# a_1235_416# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.116e+11p pd=1.34e+06u as=0p ps=0u w=360000u l=150000u
C0 vpwr VOUT 0.12fF
C1 a_1235_416# a_438_293# 0.00fF
C2 vpwr a_919_243# 0.23fF
C3 vpwr INB 0.03fF
C4 vpwr a_438_293# 0.08fF
C5 VGND a_264_22# 0.63fF
C6 VPB a_264_22# 0.16fF
C7 vpwr IN 0.01fF
C8 a_919_243# VOUT 0.00fF
C9 VGND a_1235_416# 0.00fF
C10 a_1235_416# VPB 0.00fF
C11 VOUT INB 0.00fF
C12 VOUT a_438_293# 0.01fF
C13 a_919_243# INB 0.13fF
C14 VGND vpwr 0.31fF
C15 vpwr VPB 0.35fF
C16 a_919_243# a_438_293# 0.01fF
C17 VOUT IN 0.01fF
C18 a_919_243# IN 0.03fF
C19 INB IN 0.01fF
C20 IN a_438_293# 0.03fF
C21 a_1235_416# a_264_22# 0.00fF
C22 VGND VOUT 0.05fF
C23 VOUT VPB 0.06fF
C24 VGND a_919_243# 0.59fF
C25 vpwr a_264_22# 0.14fF
C26 a_919_243# VPB 0.18fF
C27 VGND INB 0.05fF
C28 INB VPB 0.05fF
C29 VGND a_438_293# 0.01fF
C30 VPB a_438_293# 0.06fF
C31 vpwr a_1235_416# 0.00fF
C32 VGND IN 0.05fF
C33 IN VPB 0.03fF
C34 VOUT a_264_22# 0.11fF
C35 a_919_243# a_264_22# 0.28fF
C36 INB a_264_22# 0.01fF
C37 a_1235_416# VOUT 0.00fF
C38 VGND VPB 0.10fF
C39 a_438_293# a_264_22# 0.27fF
C40 a_919_243# a_1235_416# 0.00fF
C41 IN a_264_22# 0.19fF
C42 VPB VNB 2.74fF
C43 IN VNB 0.57fF
C44 INB VNB 0.62fF
C45 VOUT VNB 0.11fF
C46 a_919_243# VNB 0.26fF
C47 a_264_22# VNB 0.32fF
C48 a_438_293# VNB 0.15fF
C49 VGND VNB 1.58fF
C50 vpwr VNB 1.34fF
.ends

.subckt sky130_fd_sc_hd__o211a_1 C1 B1 A2 A1 X VGND VPWR VNB a_297_297# VPB a_510_47#
+ a_215_47# a_79_21#
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=3.8025e+11p pd=3.77e+06u as=4.55e+11p ps=4e+06u w=650000u l=150000u
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=2.275e+11p pd=2e+06u as=0p ps=0u w=650000u l=150000u
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=7.4e+11p pd=5.48e+06u as=8.7e+11p ps=7.74e+06u w=1e+06u l=150000u
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.25e+11p ps=2.65e+06u w=1e+06u l=150000u
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.9e+06u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 VGND A2 0.01fF
C1 a_297_297# VGND 0.00fF
C2 a_215_47# C1 0.00fF
C3 B1 C1 0.05fF
C4 A1 X 0.00fF
C5 VPWR A2 0.01fF
C6 a_297_297# VPWR 0.00fF
C7 a_215_47# VGND 0.20fF
C8 B1 VGND 0.01fF
C9 a_215_47# VPWR 0.01fF
C10 a_510_47# X 0.00fF
C11 B1 VPWR 0.01fF
C12 a_215_47# A2 0.04fF
C13 B1 A2 0.06fF
C14 a_297_297# a_215_47# 0.00fF
C15 a_79_21# VPB 0.03fF
C16 B1 a_215_47# 0.00fF
C17 a_79_21# X 0.03fF
C18 VPB C1 0.02fF
C19 a_79_21# A1 0.09fF
C20 VPB VGND 0.02fF
C21 X C1 0.00fF
C22 VPB VPWR 0.08fF
C23 a_79_21# a_510_47# 0.00fF
C24 X VGND 0.09fF
C25 X VPWR 0.11fF
C26 VPB A2 0.01fF
C27 A1 C1 0.00fF
C28 X A2 0.00fF
C29 VPB a_215_47# 0.00fF
C30 a_297_297# X 0.00fF
C31 B1 VPB 0.01fF
C32 A1 VGND 0.01fF
C33 A1 VPWR 0.01fF
C34 X a_215_47# 0.00fF
C35 B1 X 0.00fF
C36 a_510_47# VGND 0.00fF
C37 A1 A2 0.07fF
C38 A1 a_297_297# 0.00fF
C39 a_510_47# VPWR 0.00fF
C40 a_79_21# C1 0.07fF
C41 A1 a_215_47# 0.05fF
C42 B1 A1 0.00fF
C43 a_79_21# VGND 0.10fF
C44 a_510_47# a_215_47# 0.00fF
C45 a_79_21# VPWR 0.33fF
C46 B1 a_510_47# 0.00fF
C47 a_79_21# A2 0.04fF
C48 a_79_21# a_297_297# 0.00fF
C49 C1 VGND 0.01fF
C50 VPB X 0.01fF
C51 a_79_21# a_215_47# 0.04fF
C52 B1 a_79_21# 0.06fF
C53 VPWR C1 0.01fF
C54 VPWR VGND 0.09fF
C55 C1 A2 0.00fF
C56 A1 VPB 0.01fF
C57 VGND VNB 0.45fF
C58 VPWR VNB 0.40fF
C59 X VNB 0.10fF
C60 C1 VNB 0.18fF
C61 B1 VNB 0.08fF
C62 A2 VNB 0.09fF
C63 A1 VNB 0.08fF
C64 VPB VNB 0.78fF
C65 a_215_47# VNB 0.01fF
C66 a_79_21# VNB 0.26fF
.ends

.subckt sky130_fd_sc_hd__conb_1 LO HI VNB VPB VGND VPWR
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
C0 HI VPWR 0.07fF
C1 LO VPB 0.01fF
C2 LO VGND 0.06fF
C3 LO HI 0.07fF
C4 VGND VPB 0.02fF
C5 LO VPWR 0.21fF
C6 HI VPB 0.01fF
C7 HI VGND 0.13fF
C8 VPWR VPB 0.04fF
C9 VPWR VGND 0.04fF
C10 VGND VNB 0.38fF
C11 LO VNB 0.20fF
C12 HI VNB 0.23fF
C13 VPWR VNB 0.34fF
C14 VPB VNB 0.34fF
.ends

.subckt sky130_fd_sc_hd__mux4_2 X S0 A2 A3 S1 A1 A0 VGND VPWR VNB VPB a_193_369# a_372_413#
+ a_1281_47# a_193_47# a_1064_47# a_1060_369# a_288_47# a_397_47# a_872_316# a_1279_413#
+ a_788_316# a_600_345# a_27_47#
X0 a_600_345# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=1.16e+12p ps=1.079e+07u w=640000u l=150000u
X1 a_788_316# S1 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=1.155e+11p pd=1.39e+06u as=2.514e+11p ps=2.87e+06u w=420000u l=150000u
X2 VPWR A3 a_372_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=3.29e+11p ps=2.66e+06u w=640000u l=150000u
X3 a_872_316# a_600_345# a_788_316# VNB sky130_fd_pr__nfet_01v8 ad=2.532e+11p pd=2.88e+06u as=0p ps=0u w=420000u l=150000u
X4 VPWR S0 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X5 a_1279_413# S0 a_872_316# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.107e+11p pd=1.99e+06u as=2.538e+11p ps=2.98e+06u w=420000u l=150000u
X6 VGND a_788_316# X VNB sky130_fd_pr__nfet_01v8 ad=8.209e+11p pd=8.35e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X7 a_1060_369# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.755e+11p pd=2.33e+06u as=0p ps=0u w=640000u l=150000u
X8 a_872_316# a_27_47# a_1060_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_1281_47# a_27_47# a_872_316# VNB sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=360000u l=150000u
X10 a_193_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X11 a_1064_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.572e+11p pd=1.61e+06u as=0p ps=0u w=420000u l=150000u
X12 a_872_316# S1 a_788_316# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.458e+11p ps=1.62e+06u w=540000u l=150000u
X13 a_872_316# S0 a_1064_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 X a_788_316# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_788_316# a_600_345# a_288_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.538e+11p ps=2.98e+06u w=540000u l=150000u
X16 a_372_413# a_27_47# a_288_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND A3 a_397_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.341e+11p ps=1.5e+06u w=420000u l=150000u
X18 a_600_345# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X19 a_193_369# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.915e+11p pd=1.93e+06u as=0p ps=0u w=640000u l=150000u
X20 VPWR a_788_316# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X21 a_288_47# S0 a_193_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 a_397_47# S0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23 VGND A0 a_1281_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_288_47# a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X25 X a_788_316# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND S0 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X27 VPWR A0 a_1279_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
C0 A3 a_600_345# 0.00fF
C1 a_288_47# a_600_345# 0.13fF
C2 a_193_369# S0 0.00fF
C3 a_1279_413# S0 0.00fF
C4 VPB a_872_316# 0.02fF
C5 A2 VPWR 0.01fF
C6 a_1281_47# A0 0.00fF
C7 A1 a_872_316# 0.15fF
C8 a_1064_47# A0 0.00fF
C9 S1 VPB 0.05fF
C10 a_788_316# a_193_369# 0.00fF
C11 A0 X 0.01fF
C12 A1 S1 0.01fF
C13 a_1060_369# S0 0.00fF
C14 a_27_47# a_1281_47# 0.00fF
C15 a_788_316# a_1279_413# 0.01fF
C16 a_27_47# a_1064_47# 0.00fF
C17 VGND a_193_47# 0.00fF
C18 a_27_47# X 0.00fF
C19 a_788_316# a_1060_369# 0.00fF
C20 a_193_369# A2 0.00fF
C21 VGND a_397_47# 0.00fF
C22 A0 a_600_345# 0.00fF
C23 a_193_47# VPWR 0.00fF
C24 A3 VGND 0.03fF
C25 a_372_413# S0 0.00fF
C26 S1 a_872_316# 0.00fF
C27 a_288_47# VGND 0.08fF
C28 X VPB 0.00fF
C29 a_27_47# a_600_345# 0.01fF
C30 A1 X 0.00fF
C31 a_788_316# S0 0.06fF
C32 a_788_316# a_372_413# 0.00fF
C33 a_397_47# VPWR 0.00fF
C34 A2 S0 0.14fF
C35 A3 VPWR 0.01fF
C36 a_288_47# VPWR 0.31fF
C37 VPB a_600_345# 0.02fF
C38 A1 a_600_345# 0.02fF
C39 a_1281_47# a_872_316# 0.00fF
C40 a_1064_47# a_872_316# 0.01fF
C41 a_788_316# A2 0.00fF
C42 X a_872_316# 0.00fF
C43 S1 X 0.00fF
C44 A0 VGND 0.06fF
C45 a_193_369# a_288_47# 0.00fF
C46 a_288_47# a_1279_413# 0.00fF
C47 a_27_47# VGND 0.07fF
C48 a_193_47# S0 0.00fF
C49 a_288_47# a_1060_369# 0.00fF
C50 a_600_345# a_872_316# 0.00fF
C51 A0 VPWR 0.01fF
C52 S1 a_600_345# 0.21fF
C53 a_788_316# a_193_47# 0.00fF
C54 a_1281_47# X 0.00fF
C55 a_397_47# S0 0.00fF
C56 a_1064_47# X 0.00fF
C57 a_27_47# VPWR 0.17fF
C58 VGND VPB 0.06fF
C59 A1 VGND 0.04fF
C60 A2 a_193_47# 0.00fF
C61 A3 S0 0.05fF
C62 a_288_47# S0 0.02fF
C63 a_788_316# a_397_47# 0.00fF
C64 A3 a_372_413# 0.00fF
C65 A0 a_1279_413# 0.00fF
C66 a_288_47# a_372_413# 0.01fF
C67 a_788_316# A3 0.00fF
C68 a_193_369# a_27_47# 0.00fF
C69 a_27_47# a_1279_413# 0.00fF
C70 a_788_316# a_288_47# 0.13fF
C71 a_1281_47# a_600_345# 0.00fF
C72 a_1064_47# a_600_345# 0.00fF
C73 VPB VPWR 0.18fF
C74 A2 a_397_47# 0.00fF
C75 A1 VPWR 0.01fF
C76 X a_600_345# 0.00fF
C77 a_27_47# a_1060_369# 0.00fF
C78 A2 A3 0.00fF
C79 VGND a_872_316# 0.14fF
C80 A2 a_288_47# 0.02fF
C81 S1 VGND 0.02fF
C82 A0 S0 0.05fF
C83 a_27_47# S0 0.96fF
C84 a_872_316# VPWR 0.13fF
C85 a_27_47# a_372_413# 0.00fF
C86 a_788_316# A0 0.12fF
C87 S1 VPWR 0.03fF
C88 a_788_316# a_27_47# 0.22fF
C89 a_1281_47# VGND 0.00fF
C90 a_288_47# a_193_47# 0.00fF
C91 a_1064_47# VGND 0.00fF
C92 X VGND 0.10fF
C93 A2 A0 0.00fF
C94 a_193_369# a_872_316# 0.00fF
C95 a_872_316# a_1279_413# 0.00fF
C96 VPB S0 0.08fF
C97 A2 a_27_47# 0.10fF
C98 A3 a_397_47# 0.00fF
C99 A1 S0 0.04fF
C100 a_288_47# a_397_47# 0.00fF
C101 a_1060_369# a_872_316# 0.01fF
C102 a_788_316# VPB 0.05fF
C103 a_1281_47# VPWR 0.00fF
C104 a_1064_47# VPWR 0.00fF
C105 A3 a_288_47# 0.05fF
C106 a_788_316# A1 0.00fF
C107 X VPWR 0.14fF
C108 VGND a_600_345# 0.06fF
C109 A2 VPB 0.01fF
C110 A0 a_193_47# 0.00fF
C111 A2 A1 0.00fF
C112 a_872_316# S0 0.03fF
C113 a_27_47# a_193_47# 0.00fF
C114 a_193_369# X 0.00fF
C115 X a_1279_413# 0.00fF
C116 S1 S0 0.01fF
C117 a_372_413# a_872_316# 0.00fF
C118 a_600_345# VPWR 0.02fF
C119 A0 a_397_47# 0.00fF
C120 a_788_316# a_872_316# 0.12fF
C121 X a_1060_369# 0.00fF
C122 a_788_316# S1 0.01fF
C123 a_27_47# a_397_47# 0.00fF
C124 A3 A0 0.00fF
C125 a_288_47# A0 0.00fF
C126 A2 a_872_316# 0.00fF
C127 a_27_47# A3 0.01fF
C128 a_27_47# a_288_47# 0.36fF
C129 a_193_369# a_600_345# 0.00fF
C130 a_600_345# a_1279_413# 0.00fF
C131 A2 S1 0.00fF
C132 a_1281_47# S0 0.00fF
C133 a_1064_47# S0 0.00fF
C134 X S0 0.00fF
C135 a_1060_369# a_600_345# 0.00fF
C136 X a_372_413# 0.00fF
C137 a_788_316# a_1281_47# 0.00fF
C138 a_788_316# a_1064_47# 0.00fF
C139 A3 VPB 0.02fF
C140 a_788_316# X 0.08fF
C141 a_288_47# VPB 0.02fF
C142 VGND VPWR 0.09fF
C143 A3 A1 0.00fF
C144 a_288_47# A1 0.00fF
C145 a_193_47# a_872_316# 0.00fF
C146 A2 a_1281_47# 0.00fF
C147 A2 a_1064_47# 0.00fF
C148 a_600_345# S0 0.01fF
C149 A2 X 0.00fF
C150 a_27_47# A0 0.04fF
C151 a_600_345# a_372_413# 0.00fF
C152 a_193_369# VGND 0.00fF
C153 VGND a_1279_413# 0.00fF
C154 a_397_47# a_872_316# 0.00fF
C155 a_788_316# a_600_345# 0.01fF
C156 A3 a_872_316# 0.00fF
C157 VGND a_1060_369# 0.00fF
C158 a_288_47# a_872_316# 0.00fF
C159 A3 S1 0.13fF
C160 A2 a_600_345# 0.00fF
C161 a_288_47# S1 0.01fF
C162 A0 VPB 0.02fF
C163 A0 A1 0.00fF
C164 a_193_369# VPWR 0.00fF
C165 a_27_47# VPB 0.09fF
C166 VPWR a_1279_413# 0.00fF
C167 X a_193_47# 0.00fF
C168 a_27_47# A1 0.02fF
C169 VGND S0 0.24fF
C170 a_1060_369# VPWR 0.00fF
C171 X a_397_47# 0.00fF
C172 VGND a_372_413# 0.00fF
C173 a_288_47# a_1281_47# 0.00fF
C174 a_1064_47# a_288_47# 0.00fF
C175 a_788_316# VGND 0.07fF
C176 a_600_345# a_193_47# 0.00fF
C177 A3 X 0.00fF
C178 A0 a_872_316# 0.01fF
C179 a_288_47# X 0.00fF
C180 A1 VPB 0.03fF
C181 A0 S1 0.00fF
C182 a_27_47# a_872_316# 0.19fF
C183 VPWR S0 0.10fF
C184 A2 VGND 0.03fF
C185 a_27_47# S1 0.00fF
C186 a_372_413# VPWR 0.00fF
C187 a_600_345# a_397_47# 0.00fF
C188 a_788_316# VPWR 0.44fF
C189 X VNB 0.03fF
C190 VGND VNB 0.98fF
C191 A0 VNB 0.11fF
C192 A1 VNB 0.11fF
C193 S1 VNB 0.27fF
C194 A3 VNB 0.09fF
C195 VPWR VNB 0.86fF
C196 A2 VNB 0.08fF
C197 S0 VNB 0.46fF
C198 VPB VNB 1.67fF
C199 a_872_316# VNB 0.04fF
C200 a_600_345# VNB 0.10fF
C201 a_788_316# VNB 0.23fF
C202 a_288_47# VNB 0.03fF
C203 a_27_47# VNB 0.28fF
.ends

.subckt sky130_fd_sc_hd__nand2_1 Y B A VGND VPWR VNB VPB a_113_47#
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=5.2e+11p pd=5.04e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 Y a_113_47# 0.01fF
C1 B VPWR 0.03fF
C2 A VGND 0.01fF
C3 VPB VPWR 0.04fF
C4 VGND a_113_47# 0.00fF
C5 B A 0.05fF
C6 VPB A 0.02fF
C7 Y VGND 0.11fF
C8 VPWR A 0.03fF
C9 Y B 0.02fF
C10 VPWR a_113_47# 0.00fF
C11 Y VPB 0.00fF
C12 B VGND 0.03fF
C13 VPB VGND 0.01fF
C14 Y VPWR 0.20fF
C15 B VPB 0.02fF
C16 VPWR VGND 0.04fF
C17 Y A 0.07fF
C18 VGND VNB 0.24fF
C19 Y VNB 0.06fF
C20 VPWR VNB 0.27fF
C21 A VNB 0.15fF
C22 B VNB 0.15fF
C23 VPB VNB 0.34fF
.ends

.subckt sky130_fd_sc_hd__or2_2 B X A VPWR VGND a_39_297# VNB VPB a_121_297#
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=4.917e+11p ps=5.19e+06u w=650000u l=150000u
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=5.715e+11p pd=5.23e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 A B 0.08fF
C1 VGND A 0.03fF
C2 VPB VPWR 0.06fF
C3 a_121_297# VPWR 0.00fF
C4 VGND B 0.02fF
C5 a_39_297# A 0.17fF
C6 X A 0.01fF
C7 a_39_297# B 0.06fF
C8 VGND a_39_297# 0.10fF
C9 X B 0.00fF
C10 X VGND 0.09fF
C11 VPWR A 0.00fF
C12 VPWR B 0.01fF
C13 X a_39_297# 0.09fF
C14 VPWR VGND 0.06fF
C15 VPB A 0.01fF
C16 VPB B 0.02fF
C17 VPB VGND 0.02fF
C18 a_121_297# VGND 0.00fF
C19 VPWR a_39_297# 0.07fF
C20 X VPWR 0.13fF
C21 VPB a_39_297# 0.03fF
C22 X VPB 0.01fF
C23 a_121_297# a_39_297# 0.00fF
C24 a_121_297# X 0.00fF
C25 VGND VNB 0.33fF
C26 X VNB 0.08fF
C27 A VNB 0.10fF
C28 B VNB 0.18fF
C29 VPWR VNB 0.30fF
C30 VPB VNB 0.52fF
C31 a_39_297# VNB 0.25fF
.ends

.subckt sky130_fd_sc_hd__o311a_1 X A1 A2 A3 B1 C1 VGND VPWR VNB VPB a_368_297# a_266_47#
+ a_266_297# a_81_21# a_585_47#
X0 a_585_47# B1 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.72e+06u as=4.7125e+11p ps=4.05e+06u w=650000u l=150000u
X1 VGND A2 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=6.7925e+11p pd=4.69e+06u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=9.25e+11p pd=5.85e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3 a_81_21# C1 a_585_47# VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X5 a_266_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.6e+11p pd=2.72e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_368_297# A2 a_266_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.2e+11p pd=2.84e+06u as=0p ps=0u w=1e+06u l=150000u
X7 a_266_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_266_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_81_21# A3 a_368_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.35e+11p pd=5.07e+06u as=0p ps=0u w=1e+06u l=150000u
X10 a_81_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_81_21# a_266_47# 0.04fF
C1 X VGND 0.07fF
C2 A3 C1 0.00fF
C3 A2 A1 0.07fF
C4 VPWR C1 0.01fF
C5 VPB X 0.01fF
C6 A3 a_266_47# 0.04fF
C7 a_585_47# VGND 0.00fF
C8 a_81_21# B1 0.07fF
C9 VPWR a_266_47# 0.00fF
C10 A2 C1 0.00fF
C11 a_81_21# VGND 0.10fF
C12 X a_266_297# 0.00fF
C13 A2 a_266_47# 0.05fF
C14 a_368_297# X 0.00fF
C15 A1 C1 0.00fF
C16 A3 B1 0.08fF
C17 VPB a_81_21# 0.03fF
C18 VPWR B1 0.01fF
C19 A3 VGND 0.01fF
C20 A1 a_266_47# 0.00fF
C21 VPWR VGND 0.09fF
C22 A2 B1 0.00fF
C23 X a_585_47# 0.00fF
C24 VPB A3 0.01fF
C25 a_81_21# a_266_297# 0.01fF
C26 VPB VPWR 0.07fF
C27 a_368_297# a_81_21# 0.01fF
C28 A2 VGND 0.01fF
C29 C1 a_266_47# 0.00fF
C30 X a_81_21# 0.06fF
C31 A1 B1 0.00fF
C32 VPB A2 0.01fF
C33 A3 a_266_297# 0.00fF
C34 VPWR a_266_297# 0.00fF
C35 a_368_297# A3 0.01fF
C36 A1 VGND 0.03fF
C37 a_368_297# VPWR 0.00fF
C38 a_81_21# a_585_47# 0.00fF
C39 C1 B1 0.06fF
C40 X A3 0.00fF
C41 X VPWR 0.08fF
C42 VPB A1 0.01fF
C43 A2 a_266_297# 0.01fF
C44 a_368_297# A2 0.00fF
C45 C1 VGND 0.01fF
C46 B1 a_266_47# 0.03fF
C47 X A2 0.00fF
C48 VPWR a_585_47# 0.00fF
C49 VPB C1 0.01fF
C50 a_266_47# VGND 0.18fF
C51 a_81_21# A3 0.08fF
C52 VPWR a_81_21# 0.35fF
C53 VPB a_266_47# 0.00fF
C54 X A1 0.00fF
C55 B1 VGND 0.01fF
C56 a_81_21# A2 0.07fF
C57 X C1 0.00fF
C58 VPWR A3 0.01fF
C59 a_266_47# a_266_297# 0.00fF
C60 VPB B1 0.01fF
C61 a_368_297# a_266_47# 0.00fF
C62 X a_266_47# 0.00fF
C63 a_81_21# A1 0.12fF
C64 A3 A2 0.13fF
C65 VPB VGND 0.02fF
C66 VPWR A2 0.01fF
C67 a_266_47# a_585_47# 0.00fF
C68 a_81_21# C1 0.09fF
C69 A3 A1 0.00fF
C70 X B1 0.00fF
C71 VPWR A1 0.00fF
C72 a_266_297# VGND 0.00fF
C73 a_368_297# VGND 0.00fF
C74 VGND VNB 0.44fF
C75 VPWR VNB 0.39fF
C76 X VNB 0.10fF
C77 C1 VNB 0.15fF
C78 B1 VNB 0.08fF
C79 A3 VNB 0.09fF
C80 A2 VNB 0.08fF
C81 A1 VNB 0.08fF
C82 VPB VNB 0.78fF
C83 a_266_47# VNB 0.01fF
C84 a_81_21# VNB 0.25fF
.ends

.subckt sky130_fd_sc_hd__o221ai_1 A2 Y B1 C1 A1 B2 VGND VPWR a_213_123# VNB VPB a_109_47#
+ a_493_297# a_295_297#
X0 a_109_47# B1 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=3.409e+11p pd=3.66e+06u as=5.682e+11p ps=5.66e+06u w=650000u l=150000u
X1 Y B2 a_295_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=7.3e+11p pd=5.46e+06u as=2.4e+11p ps=2.48e+06u w=1e+06u l=150000u
X2 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.02e+12p pd=6.04e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3 a_213_123# B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_295_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_493_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A2 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X8 a_213_123# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
C0 VPWR C1 0.01fF
C1 a_493_297# A2 0.01fF
C2 a_295_297# A2 0.00fF
C3 A2 Y 0.05fF
C4 B2 B1 0.08fF
C5 VGND a_493_297# 0.00fF
C6 VGND a_295_297# 0.00fF
C7 a_213_123# B2 0.06fF
C8 VGND Y 0.03fF
C9 VPWR VPB 0.07fF
C10 a_109_47# VPWR 0.00fF
C11 a_295_297# B2 0.00fF
C12 B2 Y 0.07fF
C13 a_213_123# B1 0.03fF
C14 a_213_123# a_493_297# 0.00fF
C15 a_295_297# a_213_123# 0.00fF
C16 B1 Y 0.07fF
C17 A2 A1 0.08fF
C18 a_213_123# Y 0.02fF
C19 VGND A1 0.01fF
C20 A2 C1 0.00fF
C21 a_493_297# Y 0.00fF
C22 a_295_297# Y 0.00fF
C23 VGND C1 0.01fF
C24 B2 A1 0.00fF
C25 A2 VPB 0.01fF
C26 VGND VPB 0.02fF
C27 a_109_47# A2 0.00fF
C28 B2 C1 0.00fF
C29 a_109_47# VGND 0.09fF
C30 B1 A1 0.00fF
C31 a_213_123# A1 0.04fF
C32 B2 VPB 0.01fF
C33 a_109_47# B2 0.00fF
C34 B1 C1 0.02fF
C35 a_213_123# C1 0.00fF
C36 Y A1 0.00fF
C37 VPWR A2 0.09fF
C38 VPWR VGND 0.07fF
C39 B1 VPB 0.01fF
C40 a_213_123# VPB 0.00fF
C41 a_109_47# B1 0.00fF
C42 a_109_47# a_213_123# 0.08fF
C43 Y C1 0.09fF
C44 VPWR B2 0.01fF
C45 Y VPB 0.01fF
C46 a_109_47# a_295_297# 0.00fF
C47 a_109_47# Y 0.05fF
C48 VPWR B1 0.01fF
C49 VPWR a_213_123# 0.01fF
C50 A1 C1 0.00fF
C51 VPWR a_493_297# 0.00fF
C52 VPWR a_295_297# 0.00fF
C53 VPWR Y 0.24fF
C54 VGND A2 0.01fF
C55 A1 VPB 0.02fF
C56 a_109_47# A1 0.00fF
C57 A2 B2 0.06fF
C58 C1 VPB 0.01fF
C59 VGND B2 0.01fF
C60 a_109_47# C1 0.00fF
C61 a_109_47# VPB 0.00fF
C62 A2 B1 0.00fF
C63 a_213_123# A2 0.04fF
C64 VPWR A1 0.03fF
C65 VGND B1 0.01fF
C66 VGND a_213_123# 0.13fF
C67 VGND VNB 0.39fF
C68 VPWR VNB 0.39fF
C69 Y VNB 0.10fF
C70 A1 VNB 0.15fF
C71 A2 VNB 0.08fF
C72 B2 VNB 0.08fF
C73 B1 VNB 0.09fF
C74 C1 VNB 0.14fF
C75 VPB VNB 0.69fF
C76 a_213_123# VNB 0.04fF
C77 a_109_47# VNB 0.01fF
.ends

.subckt tempsenseInst_error CLK_REF DONE DOUT[0] DOUT[10] DOUT[11] DOUT[13] DOUT[17]
+ DOUT[18] DOUT[20] DOUT[21] DOUT[2] DOUT[3] DOUT[4] DOUT[5] DOUT[6] DOUT[7] DOUT[8]
+ RESET_COUNTERn SEL_CONV_TIME[2] SEL_CONV_TIME[3] en out DOUT[12] DOUT[14] DOUT[15]
+ DOUT[16] DOUT[19] DOUT[1] DOUT[22] DOUT[23] DOUT[9] SEL_CONV_TIME[0] SEL_CONV_TIME[1]
+ VIN VSS lc_out outb VDD
XHEADER_1 VIN VDD HEADER_1/a_508_138# VSS VSS VDD VDD HEADER
Xsky130_fd_sc_hd__decap_4_90 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__or3_1_0 SEL_CONV_TIME[1] sky130_fd_sc_hd__or3_1_0/X SEL_CONV_TIME[0]
+ sky130_fd_sc_hd__or3_1_0/C VDD VSS sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__or3_1_0/a_183_297#
+ VSS VDD sky130_fd_sc_hd__or3_1_0/a_111_297# sky130_fd_sc_hd__or3_1
Xsky130_fd_sc_hd__inv_1_4 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__inv_1_4/A VSS
+ VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__nor3_1_6 sky130_fd_sc_hd__nor3_2_3/C DOUT[11] sky130_fd_sc_hd__inv_1_8/Y
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_6/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__inv_1_48 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__inv_1_48/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_26 sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__inv_1_26/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_15 sky130_fd_sc_hd__nor3_1_0/A sky130_fd_sc_hd__inv_1_15/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_37 sky130_fd_sc_hd__nor3_2_2/A sky130_fd_sc_hd__inv_1_37/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__nor3_1_20 sky130_fd_sc_hd__nor3_2_3/C DOUT[14] sky130_fd_sc_hd__inv_1_39/Y
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_20/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_20/a_109_297# sky130_fd_sc_hd__nor3_1
XHEADER_2 VIN VDD HEADER_2/a_508_138# VSS VSS VDD VDD HEADER
Xsky130_fd_sc_hd__decap_4_91 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_80 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nor3_1_7 sky130_fd_sc_hd__nor3_2_3/C DOUT[19] sky130_fd_sc_hd__inv_1_2/Y
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_7/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__inv_1_5 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__inv_1_5/A VSS
+ VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_49 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__inv_1_49/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_27 sky130_fd_sc_hd__inv_1_27/Y sky130_fd_sc_hd__inv_1_27/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_38 sky130_fd_sc_hd__inv_1_38/Y sky130_fd_sc_hd__inv_1_38/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_16 sky130_fd_sc_hd__inv_1_17/A sky130_fd_sc_hd__inv_1_18/Y
+ VSS VIN VSS VIN sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__nor3_1_10 sky130_fd_sc_hd__nor3_2_3/C DOUT[7] sky130_fd_sc_hd__inv_1_6/Y
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_10/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_10/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__decap_4_92 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_81 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nor3_1_8 sky130_fd_sc_hd__nor3_2_3/C DOUT[6] sky130_fd_sc_hd__inv_1_3/Y
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_8/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__inv_1_6 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__inv_1_6/A VSS
+ VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_28 sky130_fd_sc_hd__inv_1_28/Y sky130_fd_sc_hd__inv_1_28/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_17 sky130_fd_sc_hd__inv_1_23/A sky130_fd_sc_hd__inv_1_17/A
+ VSS VIN VSS VIN sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_39 sky130_fd_sc_hd__inv_1_39/Y sky130_fd_sc_hd__inv_1_39/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__nor3_1_11 sky130_fd_sc_hd__nor3_2_3/C DOUT[8] sky130_fd_sc_hd__inv_1_4/Y
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_11/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_11/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__decap_4_60 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_71 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_82 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_1_7 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__inv_1_7/A VSS
+ VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__nor3_1_9 sky130_fd_sc_hd__nor3_2_3/C DOUT[3] sky130_fd_sc_hd__inv_1_5/Y
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_9/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__inv_1_29 sky130_fd_sc_hd__inv_1_29/Y sky130_fd_sc_hd__inv_1_29/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_18 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_1_21/Y
+ VSS VIN VSS VIN sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__nor3_1_12 sky130_fd_sc_hd__nor3_2_3/C DOUT[12] sky130_fd_sc_hd__inv_1_9/Y
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_12/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_12/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__dfrtp_1_0 sky130_fd_sc_hd__inv_1_26/A RESET_COUNTERn sky130_fd_sc_hd__nor3_2_1/A
+ sky130_fd_sc_hd__o211a_1_0/X VSS VDD sky130_fd_sc_hd__dfrtp_1_0/a_1462_47# sky130_fd_sc_hd__dfrtp_1_0/a_543_47#
+ VSS VDD sky130_fd_sc_hd__dfrtp_1_0/a_651_413# sky130_fd_sc_hd__dfrtp_1_0/a_193_47#
+ sky130_fd_sc_hd__dfrtp_1_0/a_805_47# sky130_fd_sc_hd__dfrtp_1_0/a_448_47# sky130_fd_sc_hd__dfrtp_1_0/a_639_47#
+ sky130_fd_sc_hd__dfrtp_1_0/a_1283_21# sky130_fd_sc_hd__dfrtp_1_0/a_761_289# sky130_fd_sc_hd__dfrtp_1_0/a_1108_47#
+ sky130_fd_sc_hd__dfrtp_1_0/a_1217_47# sky130_fd_sc_hd__dfrtp_1_0/a_1270_413# sky130_fd_sc_hd__dfrtp_1_0/a_27_47#
+ sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__a221oi_4_0 sky130_fd_sc_hd__o2111a_2_0/X sky130_fd_sc_hd__nor3_2_3/C
+ SEL_CONV_TIME[2] sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__inv_1_41/Y sky130_fd_sc_hd__mux4_2_0/X
+ VDD VSS sky130_fd_sc_hd__a221oi_4_0/a_1241_47# VSS VDD sky130_fd_sc_hd__a221oi_4_0/a_453_47#
+ sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__a221oi_4
Xsky130_fd_sc_hd__decap_4_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_61 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_50 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_83 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_1_8 sky130_fd_sc_hd__inv_1_8/Y sky130_fd_sc_hd__inv_1_8/A VSS
+ VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_19 sky130_fd_sc_hd__inv_1_22/A sky130_fd_sc_hd__inv_1_19/A
+ VSS VIN VSS VIN sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__nor3_1_13 sky130_fd_sc_hd__nor3_2_3/C DOUT[21] sky130_fd_sc_hd__inv_1_11/Y
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_13/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_13/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__dfrtp_1_1 sky130_fd_sc_hd__or2_2_0/B RESET_COUNTERn sky130_fd_sc_hd__dfrtp_1_1/D
+ CLK_REF VSS VDD sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# sky130_fd_sc_hd__dfrtp_1_1/a_543_47#
+ VSS VDD sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__dfrtp_1_1/a_193_47#
+ sky130_fd_sc_hd__dfrtp_1_1/a_805_47# sky130_fd_sc_hd__dfrtp_1_1/a_448_47# sky130_fd_sc_hd__dfrtp_1_1/a_639_47#
+ sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__dfrtp_1_1/a_1108_47#
+ sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# sky130_fd_sc_hd__dfrtp_1_1/a_27_47#
+ sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__decap_4_73 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_95 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_62 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_40 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_51 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_84 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__inv_1_9 sky130_fd_sc_hd__inv_1_9/Y sky130_fd_sc_hd__inv_1_9/A VSS
+ VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__nor2_1_0 sky130_fd_sc_hd__nor3_2_3/C DONE sky130_fd_sc_hd__nor3_2_3/B
+ VSS VDD VSS VDD sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor3_1_14 sky130_fd_sc_hd__nor3_2_3/C DOUT[10] sky130_fd_sc_hd__inv_1_13/Y
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_14/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_14/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__dfrtp_1_2 sky130_fd_sc_hd__inv_1_29/A RESET_COUNTERn sky130_fd_sc_hd__inv_1_29/Y
+ sky130_fd_sc_hd__o211a_1_1/X VSS VDD sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# sky130_fd_sc_hd__dfrtp_1_2/a_543_47#
+ VSS VDD sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__dfrtp_1_2/a_193_47#
+ sky130_fd_sc_hd__dfrtp_1_2/a_805_47# sky130_fd_sc_hd__dfrtp_1_2/a_448_47# sky130_fd_sc_hd__dfrtp_1_2/a_639_47#
+ sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__dfrtp_1_2/a_1108_47#
+ sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# sky130_fd_sc_hd__dfrtp_1_2/a_27_47#
+ sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__decap_4_96 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_74 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_41 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_52 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_30 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nor3_1_15 sky130_fd_sc_hd__nor3_2_3/C DOUT[13] sky130_fd_sc_hd__inv_1_36/Y
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_15/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_15/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__dfrtp_1_3 sky130_fd_sc_hd__or2_2_0/A RESET_COUNTERn sky130_fd_sc_hd__or2_2_0/X
+ CLK_REF VSS VDD sky130_fd_sc_hd__dfrtp_1_3/a_1462_47# sky130_fd_sc_hd__dfrtp_1_3/a_543_47#
+ VSS VDD sky130_fd_sc_hd__dfrtp_1_3/a_651_413# sky130_fd_sc_hd__dfrtp_1_3/a_193_47#
+ sky130_fd_sc_hd__dfrtp_1_3/a_805_47# sky130_fd_sc_hd__dfrtp_1_3/a_448_47# sky130_fd_sc_hd__dfrtp_1_3/a_639_47#
+ sky130_fd_sc_hd__dfrtp_1_3/a_1283_21# sky130_fd_sc_hd__dfrtp_1_3/a_761_289# sky130_fd_sc_hd__dfrtp_1_3/a_1108_47#
+ sky130_fd_sc_hd__dfrtp_1_3/a_1217_47# sky130_fd_sc_hd__dfrtp_1_3/a_1270_413# sky130_fd_sc_hd__dfrtp_1_3/a_27_47#
+ sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__decap_4_42 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_31 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_20 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_97 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_75 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_86 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_53 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_64 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nor3_1_16 sky130_fd_sc_hd__nor3_2_3/C DOUT[16] sky130_fd_sc_hd__inv_1_52/Y
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_16/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_16/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__decap_4_43 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_10 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_54 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_65 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_98 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_87 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nor3_1_17 sky130_fd_sc_hd__nor3_2_3/C DOUT[23] sky130_fd_sc_hd__inv_1_38/Y
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_17/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_17/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__or2b_1_0 SEL_CONV_TIME[0] SEL_CONV_TIME[1] sky130_fd_sc_hd__or2b_1_0/X
+ VSS VDD VSS VDD sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__or2b_1_0/a_219_297#
+ sky130_fd_sc_hd__or2b_1_0/a_301_297# sky130_fd_sc_hd__or2b_1
Xsky130_fd_sc_hd__decap_4_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_99 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_88 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_44 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_22 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_55 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_66 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nor3_1_18 sky130_fd_sc_hd__nor3_2_3/C DOUT[15] sky130_fd_sc_hd__inv_1_40/Y
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_18/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_18/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__decap_4_78 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_67 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_89 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_12 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_45 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_56 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__mux4_1_0 SEL_CONV_TIME[0] sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__mux4_1_0/X
+ SEL_CONV_TIME[1] sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__inv_1_43/A
+ VSS VDD sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__mux4_1_0/a_757_363#
+ sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__mux4_1_0/a_277_47# VSS VDD
+ sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__mux4_1_0/a_923_363#
+ sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__mux4_1_0/a_247_21#
+ sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__mux4_1_0/a_27_47#
+ sky130_fd_sc_hd__mux4_1
Xsky130_fd_sc_hd__nor3_1_19 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__nor3_1_19/Y
+ SEL_CONV_TIME[1] SEL_CONV_TIME[0] VSS VDD sky130_fd_sc_hd__nor3_1_19/a_193_297#
+ VSS VDD sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__nor3_2_0 sky130_fd_sc_hd__nor3_2_3/C DOUT[4] sky130_fd_sc_hd__nor3_2_0/A
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD VSS VDD sky130_fd_sc_hd__nor3_2_0/a_281_297#
+ sky130_fd_sc_hd__nor3_2_0/a_27_297# sky130_fd_sc_hd__nor3_2
Xsky130_fd_sc_hd__decap_4_13 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_24 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_68 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_46 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_57 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nor3_2_1 sky130_fd_sc_hd__nor3_2_3/C DOUT[0] sky130_fd_sc_hd__nor3_2_1/A
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD VSS VDD sky130_fd_sc_hd__nor3_2_1/a_281_297#
+ sky130_fd_sc_hd__nor3_2_1/a_27_297# sky130_fd_sc_hd__nor3_2
Xsky130_fd_sc_hd__decap_4_14 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_47 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_25 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_36 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_58 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_69 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nor3_2_2 sky130_fd_sc_hd__nor3_2_3/C DOUT[2] sky130_fd_sc_hd__nor3_2_2/A
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD VSS VDD sky130_fd_sc_hd__nor3_2_2/a_281_297#
+ sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__nor3_2
Xsky130_fd_sc_hd__decap_4_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_48 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_59 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_26 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nand3b_1_0 SEL_CONV_TIME[0] sky130_fd_sc_hd__inv_1_42/Y SEL_CONV_TIME[1]
+ sky130_fd_sc_hd__nand3b_1_0/Y VSS VDD VSS VDD sky130_fd_sc_hd__nand3b_1_0/a_53_93#
+ sky130_fd_sc_hd__nand3b_1_0/a_232_47# sky130_fd_sc_hd__nand3b_1_0/a_316_47# sky130_fd_sc_hd__nand3b_1
Xsky130_fd_sc_hd__nor3_2_3 sky130_fd_sc_hd__nor3_2_3/C DOUT[1] sky130_fd_sc_hd__nor3_2_3/A
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD VSS VDD sky130_fd_sc_hd__nor3_2_3/a_281_297#
+ sky130_fd_sc_hd__nor3_2_3/a_27_297# sky130_fd_sc_hd__nor3_2
Xsky130_fd_sc_hd__or3b_2_0 SEL_CONV_TIME[1] sky130_fd_sc_hd__or3b_2_0/B SEL_CONV_TIME[0]
+ sky130_fd_sc_hd__or3b_2_0/X VDD VSS VSS VDD sky130_fd_sc_hd__or3b_2_0/a_472_297#
+ sky130_fd_sc_hd__or3b_2_0/a_388_297# sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__or3b_2_0/a_27_47#
+ sky130_fd_sc_hd__or3b_2
Xsky130_fd_sc_hd__decap_4_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_38 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_27 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_49 VSS VIN VSS VIN sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nand3b_1_1 SEL_CONV_TIME[0] SEL_CONV_TIME[1] sky130_fd_sc_hd__inv_1_44/A
+ sky130_fd_sc_hd__nand3b_1_1/Y VSS VDD VSS VDD sky130_fd_sc_hd__nand3b_1_1/a_53_93#
+ sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__nand3b_1
Xsky130_fd_sc_hd__o2111a_2_0 SEL_CONV_TIME[3] sky130_fd_sc_hd__nand3b_1_1/Y sky130_fd_sc_hd__or2b_1_0/X
+ sky130_fd_sc_hd__inv_1_48/A sky130_fd_sc_hd__or3_1_0/X sky130_fd_sc_hd__o2111a_2_0/X
+ VSS VDD VSS sky130_fd_sc_hd__o2111a_2_0/a_386_47# VDD sky130_fd_sc_hd__o2111a_2_0/a_80_21#
+ sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__o2111a_2_0/a_458_47#
+ sky130_fd_sc_hd__o2111a_2
Xsky130_fd_sc_hd__decap_4_17 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_39 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_28 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_100 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_18 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_101 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_102 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfrtn_1_40 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__inv_1_53/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_53/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_40/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_40/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_40/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_40/a_805_47# sky130_fd_sc_hd__dfrtn_1_40/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__dfrtn_1_40/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# sky130_fd_sc_hd__dfrtn_1_40/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__decap_4_103 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfrtn_1_30 sky130_fd_sc_hd__inv_1_49/A sky130_fd_sc_hd__inv_1_50/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_50/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_30/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_30/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_30/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__dfrtn_1_30/a_805_47# sky130_fd_sc_hd__dfrtn_1_30/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_30/a_639_47# sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# sky130_fd_sc_hd__dfrtn_1_30/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# sky130_fd_sc_hd__dfrtn_1_30/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_41 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__inv_1_54/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_54/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_41/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_41/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_41/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__dfrtn_1_41/a_805_47# sky130_fd_sc_hd__dfrtn_1_41/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_41/a_639_47# sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__dfrtn_1_41/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# sky130_fd_sc_hd__dfrtn_1_41/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__decap_4_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfrtn_1_20 sky130_fd_sc_hd__inv_1_35/A sky130_fd_sc_hd__inv_1_30/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_30/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_20/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_20/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_20/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_20/a_805_47# sky130_fd_sc_hd__dfrtn_1_20/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_20/a_639_47# sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# sky130_fd_sc_hd__dfrtn_1_20/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# sky130_fd_sc_hd__dfrtn_1_20/a_1217_47# sky130_fd_sc_hd__dfrtn_1_20/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_31 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__inv_1_49/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_49/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_31/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_31/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_31/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_31/a_193_47# sky130_fd_sc_hd__dfrtn_1_31/a_805_47# sky130_fd_sc_hd__dfrtn_1_31/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_31/a_639_47# sky130_fd_sc_hd__dfrtn_1_31/a_1283_21# sky130_fd_sc_hd__dfrtn_1_31/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_31/a_1108_47# sky130_fd_sc_hd__dfrtn_1_31/a_1217_47# sky130_fd_sc_hd__dfrtn_1_31/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_42 sky130_fd_sc_hd__inv_1_25/A sky130_fd_sc_hd__inv_1_37/A
+ RESET_COUNTERn sky130_fd_sc_hd__nor3_2_2/A VSS VDD sky130_fd_sc_hd__dfrtn_1_42/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_42/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_42/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_42/a_193_47# sky130_fd_sc_hd__dfrtn_1_42/a_805_47# sky130_fd_sc_hd__dfrtn_1_42/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_42/a_639_47# sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# sky130_fd_sc_hd__dfrtn_1_42/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_42/a_1108_47# sky130_fd_sc_hd__dfrtn_1_42/a_1217_47# sky130_fd_sc_hd__dfrtn_1_42/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_42/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__decap_4_105 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XSLC_0 lc_out outb out SLC_0/a_919_243# SLC_0/a_1235_416# SLC_0/a_264_22# VSS SLC_0/a_438_293#
+ VSS VDD VDD SLC
Xsky130_fd_sc_hd__dfrtn_1_21 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__inv_1_35/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_35/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_21/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_21/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_21/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_21/a_193_47# sky130_fd_sc_hd__dfrtn_1_21/a_805_47# sky130_fd_sc_hd__dfrtn_1_21/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_21/a_639_47# sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# sky130_fd_sc_hd__dfrtn_1_21/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# sky130_fd_sc_hd__dfrtn_1_21/a_1217_47# sky130_fd_sc_hd__dfrtn_1_21/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_10 sky130_fd_sc_hd__inv_1_11/A sky130_fd_sc_hd__inv_1_10/A
+ RESET_COUNTERn sky130_fd_sc_hd__nor3_1_5/A VSS VDD sky130_fd_sc_hd__dfrtn_1_10/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_10/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_10/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_10/a_805_47# sky130_fd_sc_hd__dfrtn_1_10/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_10/a_639_47# sky130_fd_sc_hd__dfrtn_1_10/a_1283_21# sky130_fd_sc_hd__dfrtn_1_10/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# sky130_fd_sc_hd__dfrtn_1_10/a_1217_47# sky130_fd_sc_hd__dfrtn_1_10/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_32 sky130_fd_sc_hd__inv_1_9/A sky130_fd_sc_hd__inv_1_36/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_36/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_32/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_32/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_32/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_32/a_193_47# sky130_fd_sc_hd__dfrtn_1_32/a_805_47# sky130_fd_sc_hd__dfrtn_1_32/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_32/a_639_47# sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# sky130_fd_sc_hd__dfrtn_1_32/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# sky130_fd_sc_hd__dfrtn_1_32/a_1217_47# sky130_fd_sc_hd__dfrtn_1_32/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_32/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_33 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__inv_1_43/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_43/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_33/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_33/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_33/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_33/a_193_47# sky130_fd_sc_hd__dfrtn_1_33/a_805_47# sky130_fd_sc_hd__dfrtn_1_33/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_33/a_639_47# sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# sky130_fd_sc_hd__dfrtn_1_33/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_33/a_1108_47# sky130_fd_sc_hd__dfrtn_1_33/a_1217_47# sky130_fd_sc_hd__dfrtn_1_33/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_11 sky130_fd_sc_hd__inv_1_12/A sky130_fd_sc_hd__inv_1_11/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_11/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_11/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_11/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_11/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_11/a_805_47# sky130_fd_sc_hd__dfrtn_1_11/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_11/a_639_47# sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# sky130_fd_sc_hd__dfrtn_1_11/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# sky130_fd_sc_hd__dfrtn_1_11/a_1217_47# sky130_fd_sc_hd__dfrtn_1_11/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_22 sky130_fd_sc_hd__inv_1_36/A sky130_fd_sc_hd__inv_1_39/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_39/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_22/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_22/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_22/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_22/a_193_47# sky130_fd_sc_hd__dfrtn_1_22/a_805_47# sky130_fd_sc_hd__dfrtn_1_22/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_22/a_639_47# sky130_fd_sc_hd__dfrtn_1_22/a_1283_21# sky130_fd_sc_hd__dfrtn_1_22/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_22/a_1108_47# sky130_fd_sc_hd__dfrtn_1_22/a_1217_47# sky130_fd_sc_hd__dfrtn_1_22/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__o211a_1_0 lc_out sky130_fd_sc_hd__or2_2_0/B sky130_fd_sc_hd__nor3_2_3/C
+ sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__o211a_1_0/X VSS VDD VSS sky130_fd_sc_hd__o211a_1_0/a_297_297#
+ VDD sky130_fd_sc_hd__o211a_1_0/a_510_47# sky130_fd_sc_hd__o211a_1_0/a_215_47# sky130_fd_sc_hd__o211a_1_0/a_79_21#
+ sky130_fd_sc_hd__o211a_1
Xsky130_fd_sc_hd__dfrtn_1_34 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__or3b_2_0/B
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_51/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_34/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_34/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_34/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__dfrtn_1_34/a_805_47# sky130_fd_sc_hd__dfrtn_1_34/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_34/a_639_47# sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# sky130_fd_sc_hd__dfrtn_1_34/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# sky130_fd_sc_hd__dfrtn_1_34/a_1217_47# sky130_fd_sc_hd__dfrtn_1_34/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_12 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_0/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_0/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_12/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_12/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_12/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_12/a_805_47# sky130_fd_sc_hd__dfrtn_1_12/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_12/a_639_47# sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__dfrtn_1_12/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# sky130_fd_sc_hd__dfrtn_1_12/a_1217_47# sky130_fd_sc_hd__dfrtn_1_12/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_23 sky130_fd_sc_hd__inv_1_39/A sky130_fd_sc_hd__inv_1_40/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_40/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_23/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_23/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_23/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_23/a_193_47# sky130_fd_sc_hd__dfrtn_1_23/a_805_47# sky130_fd_sc_hd__dfrtn_1_23/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_23/a_639_47# sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# sky130_fd_sc_hd__dfrtn_1_23/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# sky130_fd_sc_hd__dfrtn_1_23/a_1217_47# sky130_fd_sc_hd__dfrtn_1_23/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__o211a_1_1 CLK_REF sky130_fd_sc_hd__or2_2_0/A sky130_fd_sc_hd__nor3_2_3/C
+ sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__o211a_1_1/X VSS VDD VSS sky130_fd_sc_hd__o211a_1_1/a_297_297#
+ VDD sky130_fd_sc_hd__o211a_1_1/a_510_47# sky130_fd_sc_hd__o211a_1_1/a_215_47# sky130_fd_sc_hd__o211a_1_1/a_79_21#
+ sky130_fd_sc_hd__o211a_1
Xsky130_fd_sc_hd__dfrtn_1_24 sky130_fd_sc_hd__inv_1_48/A sky130_fd_sc_hd__inv_1_44/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_44/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_24/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_24/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_24/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_24/a_805_47# sky130_fd_sc_hd__dfrtn_1_24/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_24/a_639_47# sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# sky130_fd_sc_hd__dfrtn_1_24/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# sky130_fd_sc_hd__dfrtn_1_24/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_35 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__inv_1_38/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_38/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_35/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_35/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_35/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_35/a_193_47# sky130_fd_sc_hd__dfrtn_1_35/a_805_47# sky130_fd_sc_hd__dfrtn_1_35/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_35/a_639_47# sky130_fd_sc_hd__dfrtn_1_35/a_1283_21# sky130_fd_sc_hd__dfrtn_1_35/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_35/a_1108_47# sky130_fd_sc_hd__dfrtn_1_35/a_1217_47# sky130_fd_sc_hd__dfrtn_1_35/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_13 sky130_fd_sc_hd__inv_1_13/A sky130_fd_sc_hd__inv_1_8/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_8/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_13/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_13/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_13/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__dfrtn_1_13/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__dfrtn_1_13/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# sky130_fd_sc_hd__dfrtn_1_13/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_25 sky130_fd_sc_hd__or3_1_0/C sky130_fd_sc_hd__inv_1_42/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_42/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_25/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_25/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_25/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__dfrtn_1_25/a_805_47# sky130_fd_sc_hd__dfrtn_1_25/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_25/a_639_47# sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# sky130_fd_sc_hd__dfrtn_1_25/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# sky130_fd_sc_hd__dfrtn_1_25/a_1217_47# sky130_fd_sc_hd__dfrtn_1_25/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_14 sky130_fd_sc_hd__inv_1_14/A sky130_fd_sc_hd__inv_1_1/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_1/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_14/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_14/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_14/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_14/a_193_47# sky130_fd_sc_hd__dfrtn_1_14/a_805_47# sky130_fd_sc_hd__dfrtn_1_14/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_14/a_639_47# sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# sky130_fd_sc_hd__dfrtn_1_14/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# sky130_fd_sc_hd__dfrtn_1_14/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_36 sky130_fd_sc_hd__inv_1_40/A sky130_fd_sc_hd__inv_1_52/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_52/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_36/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_36/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_36/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_36/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_805_47# sky130_fd_sc_hd__dfrtn_1_36/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_36/a_639_47# sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# sky130_fd_sc_hd__dfrtn_1_36/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# sky130_fd_sc_hd__dfrtn_1_36/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_36/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__decap_4_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_0 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__dfrtp_1_1/D
+ VSS VDD VSS VDD sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__dfrtn_1_37 sky130_fd_sc_hd__inv_1_32/A sky130_fd_sc_hd__inv_1_31/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_31/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_37/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_37/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_37/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__dfrtn_1_37/a_805_47# sky130_fd_sc_hd__dfrtn_1_37/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_37/a_639_47# sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# sky130_fd_sc_hd__dfrtn_1_37/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# sky130_fd_sc_hd__dfrtn_1_37/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_26 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__inv_1_45/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_45/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_26/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_26/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_26/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__dfrtn_1_26/a_805_47# sky130_fd_sc_hd__dfrtn_1_26/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_26/a_639_47# sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# sky130_fd_sc_hd__dfrtn_1_26/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# sky130_fd_sc_hd__dfrtn_1_26/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_15 sky130_fd_sc_hd__inv_1_37/A sky130_fd_sc_hd__inv_1_5/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_5/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_15/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_15/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_15/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__dfrtn_1_15/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__dfrtn_1_15/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# sky130_fd_sc_hd__dfrtn_1_15/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__decap_4_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfrtn_1_0 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_15/A
+ RESET_COUNTERn sky130_fd_sc_hd__nor3_1_0/A VSS VDD sky130_fd_sc_hd__dfrtn_1_0/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_0/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_0/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_0/a_193_47# sky130_fd_sc_hd__dfrtn_1_0/a_805_47# sky130_fd_sc_hd__dfrtn_1_0/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_0/a_639_47# sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# sky130_fd_sc_hd__dfrtn_1_0/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# sky130_fd_sc_hd__dfrtn_1_0/a_1217_47# sky130_fd_sc_hd__dfrtn_1_0/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_38 sky130_fd_sc_hd__inv_1_53/A sky130_fd_sc_hd__inv_1_27/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_27/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_38/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_38/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_38/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_38/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_805_47# sky130_fd_sc_hd__dfrtn_1_38/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_38/a_639_47# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# sky130_fd_sc_hd__dfrtn_1_38/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# sky130_fd_sc_hd__dfrtn_1_38/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_27 sky130_fd_sc_hd__inv_1_43/A sky130_fd_sc_hd__or3_1_0/C
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_46/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_27/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_27/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_27/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_27/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_805_47# sky130_fd_sc_hd__dfrtn_1_27/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_27/a_639_47# sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# sky130_fd_sc_hd__dfrtn_1_27/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# sky130_fd_sc_hd__dfrtn_1_27/a_1217_47# sky130_fd_sc_hd__dfrtn_1_27/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_27/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_16 sky130_fd_sc_hd__inv_1_26/A sky130_fd_sc_hd__inv_1_25/A
+ RESET_COUNTERn sky130_fd_sc_hd__nor3_2_3/A VSS VDD sky130_fd_sc_hd__dfrtn_1_16/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_16/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_16/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_16/a_193_47# sky130_fd_sc_hd__dfrtn_1_16/a_805_47# sky130_fd_sc_hd__dfrtn_1_16/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_16/a_639_47# sky130_fd_sc_hd__dfrtn_1_16/a_1283_21# sky130_fd_sc_hd__dfrtn_1_16/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_16/a_1108_47# sky130_fd_sc_hd__dfrtn_1_16/a_1217_47# sky130_fd_sc_hd__dfrtn_1_16/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_16/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__decap_4_2 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfrtn_1_1 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_3/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_3/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_1/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_1/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_1/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_1/a_805_47# sky130_fd_sc_hd__dfrtn_1_1/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__dfrtn_1_1/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# sky130_fd_sc_hd__dfrtn_1_1/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__mux4_2_0 sky130_fd_sc_hd__mux4_2_0/X SEL_CONV_TIME[1] sky130_fd_sc_hd__inv_1_32/A
+ sky130_fd_sc_hd__inv_1_53/A SEL_CONV_TIME[0] sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__inv_1_33/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__mux4_2_0/a_193_369# sky130_fd_sc_hd__mux4_2_0/a_372_413#
+ sky130_fd_sc_hd__mux4_2_0/a_1281_47# sky130_fd_sc_hd__mux4_2_0/a_193_47# sky130_fd_sc_hd__mux4_2_0/a_1064_47#
+ sky130_fd_sc_hd__mux4_2_0/a_1060_369# sky130_fd_sc_hd__mux4_2_0/a_288_47# sky130_fd_sc_hd__mux4_2_0/a_397_47#
+ sky130_fd_sc_hd__mux4_2_0/a_872_316# sky130_fd_sc_hd__mux4_2_0/a_1279_413# sky130_fd_sc_hd__mux4_2_0/a_788_316#
+ sky130_fd_sc_hd__mux4_2_0/a_600_345# sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__mux4_2
Xsky130_fd_sc_hd__nand2_1_0 sky130_fd_sc_hd__inv_1_19/A sky130_fd_sc_hd__inv_1_23/A
+ en VSS VIN VSS VIN sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__inv_1_50 sky130_fd_sc_hd__inv_1_50/Y sky130_fd_sc_hd__inv_1_50/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__dfrtn_1_39 sky130_fd_sc_hd__inv_1_33/A sky130_fd_sc_hd__inv_1_32/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_32/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_39/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_39/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_39/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_39/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_805_47# sky130_fd_sc_hd__dfrtn_1_39/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_39/a_639_47# sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# sky130_fd_sc_hd__dfrtn_1_39/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# sky130_fd_sc_hd__dfrtn_1_39/a_1217_47# sky130_fd_sc_hd__dfrtn_1_39/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_28 sky130_fd_sc_hd__inv_1_42/A sky130_fd_sc_hd__inv_1_48/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_48/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_28/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_28/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_28/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_28/a_193_47# sky130_fd_sc_hd__dfrtn_1_28/a_805_47# sky130_fd_sc_hd__dfrtn_1_28/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_28/a_639_47# sky130_fd_sc_hd__dfrtn_1_28/a_1283_21# sky130_fd_sc_hd__dfrtn_1_28/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_28/a_1108_47# sky130_fd_sc_hd__dfrtn_1_28/a_1217_47# sky130_fd_sc_hd__dfrtn_1_28/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_17 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__inv_1_28/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_28/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_17/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_17/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_17/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_17/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_805_47# sky130_fd_sc_hd__dfrtn_1_17/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_17/a_639_47# sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# sky130_fd_sc_hd__dfrtn_1_17/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# sky130_fd_sc_hd__dfrtn_1_17/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__or2_2_0 sky130_fd_sc_hd__or2_2_0/B sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__or2_2_0/A
+ VDD VSS sky130_fd_sc_hd__or2_2_0/a_39_297# VSS VDD sky130_fd_sc_hd__or2_2_0/a_121_297#
+ sky130_fd_sc_hd__or2_2
Xsky130_fd_sc_hd__decap_4_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfrtn_1_2 sky130_fd_sc_hd__inv_1_6/A sky130_fd_sc_hd__inv_1_4/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_4/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_2/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_2/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_2/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_805_47# sky130_fd_sc_hd__dfrtn_1_2/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_2/a_639_47# sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_2/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__dfrtn_1_2/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__o311a_1_0 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__inv_1_41/Y
+ sky130_fd_sc_hd__nor3_1_19/Y sky130_fd_sc_hd__o311a_1_0/A3 sky130_fd_sc_hd__nand2_1_1/Y
+ SEL_CONV_TIME[2] VSS VDD VSS VDD sky130_fd_sc_hd__o311a_1_0/a_368_297# sky130_fd_sc_hd__o311a_1_0/a_266_47#
+ sky130_fd_sc_hd__o311a_1_0/a_266_297# sky130_fd_sc_hd__o311a_1_0/a_81_21# sky130_fd_sc_hd__o311a_1_0/a_585_47#
+ sky130_fd_sc_hd__o311a_1
Xsky130_fd_sc_hd__nand2_1_1 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__mux4_1_0/X
+ sky130_fd_sc_hd__inv_1_41/Y VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1_1/a_113_47#
+ sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__inv_1_51 sky130_fd_sc_hd__inv_1_51/Y sky130_fd_sc_hd__or3b_2_0/B
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_40 sky130_fd_sc_hd__inv_1_40/Y sky130_fd_sc_hd__inv_1_40/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__dfrtn_1_29 sky130_fd_sc_hd__inv_1_44/A sky130_fd_sc_hd__inv_1_47/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_47/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_29/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_29/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_29/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__dfrtn_1_29/a_805_47# sky130_fd_sc_hd__dfrtn_1_29/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_29/a_639_47# sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# sky130_fd_sc_hd__dfrtn_1_29/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# sky130_fd_sc_hd__dfrtn_1_29/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__dfrtn_1_18 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__inv_1_33/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_33/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_18/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_18/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_18/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_18/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_805_47# sky130_fd_sc_hd__dfrtn_1_18/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_18/a_639_47# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# sky130_fd_sc_hd__dfrtn_1_18/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# sky130_fd_sc_hd__dfrtn_1_18/a_1217_47# sky130_fd_sc_hd__dfrtn_1_18/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_18/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__decap_4_4 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfrtn_1_3 sky130_fd_sc_hd__inv_1_5/A sky130_fd_sc_hd__inv_1_14/A
+ RESET_COUNTERn sky130_fd_sc_hd__nor3_2_0/A VSS VDD sky130_fd_sc_hd__dfrtn_1_3/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_3/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_3/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_3/a_805_47# sky130_fd_sc_hd__dfrtn_1_3/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_3/a_639_47# sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# sky130_fd_sc_hd__dfrtn_1_3/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# sky130_fd_sc_hd__dfrtn_1_3/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__nand2_1_2 sky130_fd_sc_hd__nand2_1_2/Y SEL_CONV_TIME[0] SEL_CONV_TIME[1]
+ VSS VDD VSS VDD sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__inv_1_30 sky130_fd_sc_hd__inv_1_30/Y sky130_fd_sc_hd__inv_1_30/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_41 sky130_fd_sc_hd__inv_1_41/Y SEL_CONV_TIME[3] VSS VDD VSS
+ VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_52 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__inv_1_52/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__dfrtn_1_19 sky130_fd_sc_hd__inv_1_28/A sky130_fd_sc_hd__inv_1_34/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_34/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_19/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_19/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_19/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_19/a_193_47# sky130_fd_sc_hd__dfrtn_1_19/a_805_47# sky130_fd_sc_hd__dfrtn_1_19/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_19/a_639_47# sky130_fd_sc_hd__dfrtn_1_19/a_1283_21# sky130_fd_sc_hd__dfrtn_1_19/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_19/a_1108_47# sky130_fd_sc_hd__dfrtn_1_19/a_1217_47# sky130_fd_sc_hd__dfrtn_1_19/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_19/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__decap_4_5 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfrtn_1_4 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_7/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_7/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_4/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_4/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_4/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_4/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_805_47# sky130_fd_sc_hd__dfrtn_1_4/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_4/a_639_47# sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# sky130_fd_sc_hd__dfrtn_1_4/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# sky130_fd_sc_hd__dfrtn_1_4/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__nor3_1_0 sky130_fd_sc_hd__nor3_2_3/C DOUT[18] sky130_fd_sc_hd__nor3_1_0/A
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_0/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_0/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__inv_1_31 sky130_fd_sc_hd__inv_1_31/Y sky130_fd_sc_hd__inv_1_31/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_53 sky130_fd_sc_hd__inv_1_53/Y sky130_fd_sc_hd__inv_1_53/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_42 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_42/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_20 out sky130_fd_sc_hd__inv_1_23/A VSS VIN VSS VIN sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_6 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfrtn_1_5 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_13/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_13/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_5/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_5/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_5/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_805_47# sky130_fd_sc_hd__dfrtn_1_5/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_5/a_639_47# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# sky130_fd_sc_hd__dfrtn_1_5/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# sky130_fd_sc_hd__dfrtn_1_5/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__nor3_1_1 sky130_fd_sc_hd__nor3_2_3/C DOUT[17] sky130_fd_sc_hd__inv_1_0/Y
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_1/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_1/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__o221ai_1_0 sky130_fd_sc_hd__or2b_1_0/X sky130_fd_sc_hd__o311a_1_0/A3
+ sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__or3b_2_0/X sky130_fd_sc_hd__inv_1_49/A
+ sky130_fd_sc_hd__inv_1_50/A VSS VDD sky130_fd_sc_hd__o221ai_1_0/a_213_123# VSS VDD
+ sky130_fd_sc_hd__o221ai_1_0/a_109_47# sky130_fd_sc_hd__o221ai_1_0/a_493_297# sky130_fd_sc_hd__o221ai_1_0/a_295_297#
+ sky130_fd_sc_hd__o221ai_1
Xsky130_fd_sc_hd__inv_1_32 sky130_fd_sc_hd__inv_1_32/Y sky130_fd_sc_hd__inv_1_32/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_10 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__inv_1_10/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_21 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__inv_1_22/Y
+ VSS VIN VSS VIN sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_43 sky130_fd_sc_hd__inv_1_43/Y sky130_fd_sc_hd__inv_1_43/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_54 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__inv_1_54/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfrtn_1_6 sky130_fd_sc_hd__inv_1_15/A sky130_fd_sc_hd__inv_1_2/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_2/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_6/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_6/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_6/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__dfrtn_1_6/a_805_47# sky130_fd_sc_hd__dfrtn_1_6/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_6/a_639_47# sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# sky130_fd_sc_hd__dfrtn_1_6/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# sky130_fd_sc_hd__dfrtn_1_6/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__nor3_1_2 sky130_fd_sc_hd__nor3_2_3/C DOUT[5] sky130_fd_sc_hd__inv_1_1/Y
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_2/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_2/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__inv_1_0 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__inv_1_0/A VSS
+ VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_44 sky130_fd_sc_hd__inv_1_44/Y sky130_fd_sc_hd__inv_1_44/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_33 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__inv_1_33/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_22 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__inv_1_22/A
+ VSS VIN VSS VIN sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_11 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__inv_1_11/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfrtn_1_7 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_6/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_6/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_7/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_7/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_7/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_7/a_193_47# sky130_fd_sc_hd__dfrtn_1_7/a_805_47# sky130_fd_sc_hd__dfrtn_1_7/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_7/a_639_47# sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# sky130_fd_sc_hd__dfrtn_1_7/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# sky130_fd_sc_hd__dfrtn_1_7/a_1217_47# sky130_fd_sc_hd__dfrtn_1_7/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_7/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__nor3_1_3 sky130_fd_sc_hd__nor3_2_3/C DOUT[9] sky130_fd_sc_hd__inv_1_7/Y
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_3/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_3/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__inv_1_1 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__inv_1_1/A VSS
+ VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_34 sky130_fd_sc_hd__inv_1_34/Y sky130_fd_sc_hd__inv_1_34/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_45 sky130_fd_sc_hd__inv_1_45/Y sky130_fd_sc_hd__inv_1_45/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_12 sky130_fd_sc_hd__nor3_1_4/A sky130_fd_sc_hd__inv_1_12/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_23 sky130_fd_sc_hd__inv_1_24/A sky130_fd_sc_hd__inv_1_23/A
+ VSS VIN VSS VIN sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__decap_4_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfrtn_1_8 sky130_fd_sc_hd__inv_1_8/A sky130_fd_sc_hd__inv_1_9/A
+ RESET_COUNTERn sky130_fd_sc_hd__inv_1_9/Y VSS VDD sky130_fd_sc_hd__dfrtn_1_8/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_8/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_8/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_8/a_193_47# sky130_fd_sc_hd__dfrtn_1_8/a_805_47# sky130_fd_sc_hd__dfrtn_1_8/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_8/a_639_47# sky130_fd_sc_hd__dfrtn_1_8/a_1283_21# sky130_fd_sc_hd__dfrtn_1_8/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_8/a_1108_47# sky130_fd_sc_hd__dfrtn_1_8/a_1217_47# sky130_fd_sc_hd__dfrtn_1_8/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_8/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__nor3_1_4 sky130_fd_sc_hd__nor3_2_3/C DOUT[20] sky130_fd_sc_hd__nor3_1_4/A
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_4/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_4/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__inv_1_2 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__inv_1_2/A VSS
+ VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_35 sky130_fd_sc_hd__inv_1_35/Y sky130_fd_sc_hd__inv_1_35/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_46 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__or3_1_0/C
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_13 sky130_fd_sc_hd__inv_1_13/Y sky130_fd_sc_hd__inv_1_13/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_24 outb sky130_fd_sc_hd__inv_1_24/A VSS VIN VSS VIN sky130_fd_sc_hd__inv_1
XHEADER_0 VIN VDD HEADER_0/a_508_138# VSS VSS VDD VDD HEADER
Xsky130_fd_sc_hd__dfrtn_1_9 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_12/A
+ RESET_COUNTERn sky130_fd_sc_hd__nor3_1_4/A VSS VDD sky130_fd_sc_hd__dfrtn_1_9/a_1462_47#
+ sky130_fd_sc_hd__dfrtn_1_9/a_543_47# VSS VDD sky130_fd_sc_hd__dfrtn_1_9/a_651_413#
+ sky130_fd_sc_hd__dfrtn_1_9/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_805_47# sky130_fd_sc_hd__dfrtn_1_9/a_448_47#
+ sky130_fd_sc_hd__dfrtn_1_9/a_639_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# sky130_fd_sc_hd__dfrtn_1_9/a_761_289#
+ sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# sky130_fd_sc_hd__dfrtn_1_9/a_1270_413#
+ sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__dfrtn_1
Xsky130_fd_sc_hd__nor3_1_5 sky130_fd_sc_hd__nor3_2_3/C DOUT[22] sky130_fd_sc_hd__nor3_1_5/A
+ sky130_fd_sc_hd__nor3_2_3/B VSS VDD sky130_fd_sc_hd__nor3_1_5/a_193_297# VSS VDD
+ sky130_fd_sc_hd__nor3_1_5/a_109_297# sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__inv_1_3 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_3/A VSS
+ VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_14 sky130_fd_sc_hd__nor3_2_0/A sky130_fd_sc_hd__inv_1_14/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_47 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__inv_1_47/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_25 sky130_fd_sc_hd__nor3_2_3/A sky130_fd_sc_hd__inv_1_25/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_36 sky130_fd_sc_hd__inv_1_36/Y sky130_fd_sc_hd__inv_1_36/A
+ VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
C0 sky130_fd_sc_hd__dfrtn_1_20/a_651_413# RESET_COUNTERn 0.01fF
C1 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# SEL_CONV_TIME[0] 0.00fF
C2 sky130_fd_sc_hd__inv_1_30/Y RESET_COUNTERn 0.04fF
C3 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C4 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__inv_1_29/Y 0.00fF
C5 DOUT[1] sky130_fd_sc_hd__dfrtn_1_23/a_805_47# 0.00fF
C6 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C7 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# 0.01fF
C8 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_18/a_761_289# 0.00fF
C9 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_18/a_543_47# 0.00fF
C10 sky130_fd_sc_hd__dfrtn_1_18/a_1270_413# DOUT[2] 0.00fF
C11 sky130_fd_sc_hd__dfrtn_1_42/a_761_289# sky130_fd_sc_hd__inv_1_25/A 0.00fF
C12 sky130_fd_sc_hd__dfrtn_1_32/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C13 sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# VDD 0.10fF
C14 sky130_fd_sc_hd__nor3_1_19/Y sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C15 sky130_fd_sc_hd__inv_1_3/A DOUT[14] 0.02fF
C16 sky130_fd_sc_hd__nand3b_1_0/a_53_93# SEL_CONV_TIME[0] 0.01fF
C17 sky130_fd_sc_hd__dfrtn_1_3/a_761_289# DOUT[11] 0.01fF
C18 sky130_fd_sc_hd__dfrtn_1_4/a_761_289# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C19 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C20 sky130_fd_sc_hd__dfrtn_1_36/a_543_47# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C21 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__nand3b_1_0/Y 0.00fF
C22 sky130_fd_sc_hd__dfrtn_1_36/a_761_289# sky130_fd_sc_hd__inv_1_52/Y 0.02fF
C23 sky130_fd_sc_hd__inv_1_44/A DOUT[21] 0.04fF
C24 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__inv_1_6/Y 0.01fF
C25 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__or2_2_0/A 0.24fF
C26 sky130_fd_sc_hd__mux4_1_0/a_1478_413# RESET_COUNTERn 0.01fF
C27 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_26/a_543_47# 0.01fF
C28 sky130_fd_sc_hd__dfrtn_1_10/a_1462_47# RESET_COUNTERn 0.00fF
C29 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# sky130_fd_sc_hd__dfrtn_1_28/a_27_47# 0.00fF
C30 sky130_fd_sc_hd__o211a_1_0/a_297_297# RESET_COUNTERn 0.00fF
C31 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.00fF
C32 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_24/a_543_47# 0.00fF
C33 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_31/a_639_47# 0.00fF
C34 sky130_fd_sc_hd__or3b_2_0/a_472_297# sky130_fd_sc_hd__dfrtn_1_31/a_448_47# 0.00fF
C35 sky130_fd_sc_hd__or3b_2_0/a_388_297# sky130_fd_sc_hd__dfrtn_1_31/a_651_413# 0.00fF
C36 sky130_fd_sc_hd__inv_1_2/Y VIN 0.18fF
C37 sky130_fd_sc_hd__dfrtn_1_17/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C38 sky130_fd_sc_hd__dfrtn_1_17/a_1462_47# VDD 0.00fF
C39 sky130_fd_sc_hd__dfrtn_1_28/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C40 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# sky130_fd_sc_hd__nor3_2_3/A 0.02fF
C41 sky130_fd_sc_hd__nor3_2_3/C DOUT[14] 0.11fF
C42 sky130_fd_sc_hd__dfrtn_1_0/a_543_47# sky130_fd_sc_hd__nor3_1_0/a_193_297# 0.00fF
C43 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# VDD 0.08fF
C44 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C45 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__inv_1_33/A 0.69fF
C46 sky130_fd_sc_hd__inv_1_15/A DOUT[18] 0.10fF
C47 sky130_fd_sc_hd__o311a_1_0/A3 sky130_fd_sc_hd__inv_1_44/A 0.07fF
C48 SEL_CONV_TIME[0] sky130_fd_sc_hd__inv_1_43/A 0.16fF
C49 sky130_fd_sc_hd__dfrtn_1_22/a_1270_413# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C50 sky130_fd_sc_hd__inv_1_7/Y DOUT[11] 0.00fF
C51 DOUT[4] sky130_fd_sc_hd__dfrtn_1_30/a_761_289# 0.00fF
C52 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# -0.00fF
C53 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# -0.00fF
C54 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_448_47# 0.00fF
C55 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C56 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.00fF
C57 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# 0.00fF
C58 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C59 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C60 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__inv_1_45/Y 0.01fF
C61 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# 0.00fF
C62 sky130_fd_sc_hd__dfrtn_1_31/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C63 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__nor3_2_3/B 0.08fF
C64 sky130_fd_sc_hd__dfrtn_1_31/a_805_47# VDD 0.00fF
C65 sky130_fd_sc_hd__mux4_2_0/a_1281_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C66 sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C67 sky130_fd_sc_hd__dfrtn_1_28/a_1108_47# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C68 sky130_fd_sc_hd__mux4_2_0/a_397_47# SEL_CONV_TIME[0] 0.00fF
C69 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C70 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C71 sky130_fd_sc_hd__dfrtn_1_35/a_639_47# RESET_COUNTERn 0.00fF
C72 sky130_fd_sc_hd__nor3_1_4/a_193_297# DOUT[14] 0.00fF
C73 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_639_47# -0.00fF
C74 sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C75 CLK_REF sky130_fd_sc_hd__dfrtn_1_21/a_805_47# 0.00fF
C76 sky130_fd_sc_hd__nor3_1_11/a_193_297# DOUT[6] 0.00fF
C77 sky130_fd_sc_hd__nor3_1_11/a_109_297# DOUT[7] 0.00fF
C78 sky130_fd_sc_hd__nand3b_1_1/Y sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C79 sky130_fd_sc_hd__dfrtn_1_29/a_805_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C80 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# DOUT[3] 0.00fF
C81 sky130_fd_sc_hd__dfrtp_1_1/a_448_47# RESET_COUNTERn -0.00fF
C82 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__inv_1_40/A 0.01fF
C83 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__inv_1_48/A 0.01fF
C84 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# 0.00fF
C85 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# 0.00fF
C86 sky130_fd_sc_hd__dfrtp_1_3/a_543_47# sky130_fd_sc_hd__dfrtn_1_17/a_761_289# 0.00fF
C87 sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# sky130_fd_sc_hd__inv_1_31/A 0.00fF
C88 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C89 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C90 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_38/a_1462_47# 0.00fF
C91 sky130_fd_sc_hd__dfrtn_1_34/a_651_413# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C92 sky130_fd_sc_hd__dfrtn_1_34/a_1270_413# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C93 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C94 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_18/a_805_47# 0.00fF
C95 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C96 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__dfrtn_1_29/a_761_289# 0.00fF
C97 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__dfrtn_1_29/a_543_47# 0.00fF
C98 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# 0.00fF
C99 sky130_fd_sc_hd__dfrtn_1_10/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C100 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# sky130_fd_sc_hd__inv_1_7/A 0.01fF
C101 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# CLK_REF 0.00fF
C102 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C103 sky130_fd_sc_hd__dfrtp_1_3/a_1283_21# VDD 0.11fF
C104 sky130_fd_sc_hd__dfrtp_1_3/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C105 VDD sky130_fd_sc_hd__o211a_1_0/X 0.22fF
C106 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# SEL_CONV_TIME[1] 0.01fF
C107 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_21/a_193_47# 0.01fF
C108 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_21/a_651_413# 0.00fF
C109 sky130_fd_sc_hd__o311a_1_0/a_266_47# RESET_COUNTERn 0.00fF
C110 sky130_fd_sc_hd__dfrtp_1_3/a_1217_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C111 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C112 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# 0.00fF
C113 sky130_fd_sc_hd__dfrtn_1_27/a_651_413# SEL_CONV_TIME[0] 0.00fF
C114 sky130_fd_sc_hd__mux4_2_0/a_1279_413# DOUT[21] 0.00fF
C115 sky130_fd_sc_hd__mux4_2_0/a_788_316# RESET_COUNTERn 0.00fF
C116 sky130_fd_sc_hd__dfrtn_1_23/a_639_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C117 sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# sky130_fd_sc_hd__dfrtn_1_28/a_639_47# 0.00fF
C118 sky130_fd_sc_hd__dfrtn_1_25/a_1462_47# sky130_fd_sc_hd__dfrtn_1_28/a_193_47# 0.00fF
C119 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_1/D 0.11fF
C120 sky130_fd_sc_hd__or2b_1_0/X sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C121 sky130_fd_sc_hd__nor3_2_2/A DOUT[2] 0.01fF
C122 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_36/a_1270_413# 0.00fF
C123 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_761_289# -0.00fF
C124 sky130_fd_sc_hd__dfrtn_1_14/a_651_413# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C125 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__o211a_1_1/X 0.00fF
C126 sky130_fd_sc_hd__dfrtn_1_42/a_1217_47# sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C127 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# RESET_COUNTERn 0.02fF
C128 sky130_fd_sc_hd__dfrtn_1_4/a_639_47# DOUT[11] 0.00fF
C129 sky130_fd_sc_hd__o211a_1_1/a_297_297# sky130_fd_sc_hd__o211a_1_1/X 0.00fF
C130 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__inv_1_35/Y 0.00fF
C131 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__dfrtn_1_33/a_448_47# -0.00fF
C132 sky130_fd_sc_hd__inv_1_10/A VDD 1.43fF
C133 sky130_fd_sc_hd__dfrtn_1_14/a_805_47# DOUT[9] 0.00fF
C134 sky130_fd_sc_hd__dfrtn_1_0/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C135 sky130_fd_sc_hd__dfrtn_1_35/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C136 sky130_fd_sc_hd__nor3_1_20/a_193_297# RESET_COUNTERn 0.00fF
C137 sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# VDD 0.00fF
C138 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C139 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# DOUT[19] 0.00fF
C140 sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C141 sky130_fd_sc_hd__mux4_1_0/a_1478_413# SEL_CONV_TIME[3] 0.00fF
C142 sky130_fd_sc_hd__dfrtn_1_41/a_1270_413# RESET_COUNTERn 0.00fF
C143 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_34/a_639_47# 0.00fF
C144 DOUT[2] sky130_fd_sc_hd__inv_1_53/A 0.26fF
C145 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C146 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# VDD 0.07fF
C147 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_7/A 0.13fF
C148 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C149 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C150 sky130_fd_sc_hd__mux4_2_0/a_1279_413# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C151 sky130_fd_sc_hd__dfrtn_1_19/a_805_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C152 sky130_fd_sc_hd__dfrtn_1_3/a_639_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C153 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.00fF
C154 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__o211a_1_1/a_215_47# 0.00fF
C155 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__o211a_1_1/a_510_47# 0.00fF
C156 sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C157 sky130_fd_sc_hd__dfrtn_1_20/a_543_47# sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.00fF
C158 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__o211a_1_1/X 0.00fF
C159 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_543_47# 0.00fF
C160 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C161 sky130_fd_sc_hd__dfrtn_1_23/a_543_47# sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C162 sky130_fd_sc_hd__dfrtn_1_27/a_193_47# RESET_COUNTERn 0.19fF
C163 sky130_fd_sc_hd__dfrtn_1_27/a_448_47# DOUT[21] 0.00fF
C164 sky130_fd_sc_hd__nor3_1_1/a_193_297# DOUT[17] -0.00fF
C165 sky130_fd_sc_hd__dfrtn_1_38/a_761_289# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C166 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C167 sky130_fd_sc_hd__dfrtn_1_35/a_761_289# sky130_fd_sc_hd__inv_1_38/A 0.01fF
C168 sky130_fd_sc_hd__dfrtn_1_3/a_651_413# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C169 sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C170 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__dfrtn_1_25/a_27_47# 0.00fF
C171 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__dfrtn_1_25/a_193_47# 0.00fF
C172 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_25/a_448_47# 0.00fF
C173 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_25/a_639_47# 0.00fF
C174 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# 0.00fF
C175 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__inv_1_4/Y 0.01fF
C176 VDD DOUT[3] 0.62fF
C177 sky130_fd_sc_hd__o311a_1_0/a_266_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C178 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# DOUT[2] 0.00fF
C179 sky130_fd_sc_hd__dfrtn_1_12/a_1462_47# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C180 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__mux4_2_0/a_872_316# 0.00fF
C181 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# sky130_fd_sc_hd__mux4_2_0/a_372_413# 0.00fF
C182 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C183 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.00fF
C184 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C185 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# sky130_fd_sc_hd__mux4_2_0/a_600_345# 0.00fF
C186 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# sky130_fd_sc_hd__mux4_2_0/a_193_369# 0.00fF
C187 DOUT[22] sky130_fd_sc_hd__inv_1_15/A 0.02fF
C188 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__inv_1_38/Y 0.01fF
C189 sky130_fd_sc_hd__inv_1_37/A sky130_fd_sc_hd__inv_1_12/A 0.18fF
C190 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C191 sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C192 sky130_fd_sc_hd__mux4_2_0/a_288_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C193 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# sky130_fd_sc_hd__nor3_1_2/a_109_297# 0.00fF
C194 sky130_fd_sc_hd__or2_2_0/a_39_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C195 sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C196 sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C197 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C198 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# 0.00fF
C199 sky130_fd_sc_hd__a221oi_4_0/a_453_47# SEL_CONV_TIME[0] 0.00fF
C200 sky130_fd_sc_hd__inv_1_2/A VDD 0.72fF
C201 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# RESET_COUNTERn 0.03fF
C202 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__inv_1_13/Y 0.02fF
C203 sky130_fd_sc_hd__nor3_1_10/a_109_297# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C204 sky130_fd_sc_hd__dfrtn_1_33/a_761_289# sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# 0.00fF
C205 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# 0.00fF
C206 VDD DOUT[5] 0.99fF
C207 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C208 sky130_fd_sc_hd__dfrtn_1_22/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C209 sky130_fd_sc_hd__dfrtn_1_4/a_543_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C210 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C211 sky130_fd_sc_hd__dfrtn_1_22/a_448_47# VDD 0.01fF
C212 DOUT[1] sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# 0.00fF
C213 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C214 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# RESET_COUNTERn 0.01fF
C215 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_761_289# -0.00fF
C216 sky130_fd_sc_hd__dfrtn_1_41/a_639_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C217 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__dfrtn_1_24/a_651_413# 0.00fF
C218 sky130_fd_sc_hd__dfrtn_1_28/a_1270_413# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C219 sky130_fd_sc_hd__dfrtn_1_41/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C220 DOUT[4] sky130_fd_sc_hd__dfrtn_1_34/a_639_47# 0.00fF
C221 sky130_fd_sc_hd__or3b_2_0/a_27_47# SEL_CONV_TIME[0] 0.02fF
C222 sky130_fd_sc_hd__inv_1_5/Y RESET_COUNTERn 0.57fF
C223 sky130_fd_sc_hd__dfrtn_1_18/a_27_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C224 sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# sky130_fd_sc_hd__dfrtp_1_1/D 0.00fF
C225 sky130_fd_sc_hd__inv_1_30/A CLK_REF 0.00fF
C226 sky130_fd_sc_hd__dfrtn_1_23/a_651_413# sky130_fd_sc_hd__inv_1_40/A 0.00fF
C227 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__inv_1_45/A 0.16fF
C228 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__dfrtp_1_1/a_761_289# 0.00fF
C229 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/a_193_47# 0.00fF
C230 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.00fF
C231 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C232 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C233 sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C234 sky130_fd_sc_hd__dfrtn_1_8/a_1283_21# sky130_fd_sc_hd__inv_1_9/A 0.01fF
C235 sky130_fd_sc_hd__o311a_1_0/a_266_47# SEL_CONV_TIME[3] 0.00fF
C236 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_10/a_639_47# 0.00fF
C237 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C238 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_543_47# 0.00fF
C239 sky130_fd_sc_hd__dfrtp_1_1/a_639_47# DOUT[23] 0.00fF
C240 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# DOUT[19] 0.00fF
C241 sky130_fd_sc_hd__dfrtn_1_8/a_639_47# DOUT[12] 0.00fF
C242 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C243 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C244 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__inv_1_12/A 0.01fF
C245 sky130_fd_sc_hd__mux4_2_0/a_788_316# SEL_CONV_TIME[3] 0.01fF
C246 sky130_fd_sc_hd__nor3_2_1/A SLC_0/a_438_293# 0.00fF
C247 sky130_fd_sc_hd__dfrtn_1_16/a_1283_21# VDD 0.10fF
C248 sky130_fd_sc_hd__dfrtn_1_16/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C249 sky130_fd_sc_hd__dfrtn_1_8/a_27_47# VDD 0.19fF
C250 sky130_fd_sc_hd__dfrtn_1_40/a_1270_413# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C251 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_651_413# -0.00fF
C252 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C253 sky130_fd_sc_hd__a221oi_4_0/a_471_297# DOUT[21] 0.00fF
C254 sky130_fd_sc_hd__nor3_2_3/C SEL_CONV_TIME[0] 0.05fF
C255 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__inv_1_8/Y 0.01fF
C256 HEADER_2/a_508_138# HEADER_1/a_508_138# 0.00fF
C257 CLK_REF sky130_fd_sc_hd__dfrtn_1_19/a_639_47# 0.00fF
C258 sky130_fd_sc_hd__nor3_2_2/a_281_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C259 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_20/a_761_289# 0.01fF
C260 sky130_fd_sc_hd__dfrtn_1_20/a_1462_47# sky130_fd_sc_hd__dfrtn_1_18/a_543_47# 0.00fF
C261 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C262 sky130_fd_sc_hd__dfrtn_1_18/a_1270_413# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C263 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# SEL_CONV_TIME[0] 0.02fF
C264 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# sky130_fd_sc_hd__nor3_2_1/A 0.01fF
C265 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C266 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_34/a_639_47# 0.00fF
C267 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_40/a_543_47# -0.00fF
C268 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# DOUT[2] 0.00fF
C269 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# sky130_fd_sc_hd__o211a_1_0/a_215_47# 0.00fF
C270 sky130_fd_sc_hd__dfrtn_1_23/a_1462_47# sky130_fd_sc_hd__dfrtn_1_36/a_543_47# 0.00fF
C271 sky130_fd_sc_hd__dfrtn_1_23/a_1270_413# sky130_fd_sc_hd__dfrtn_1_36/a_651_413# 0.00fF
C272 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C273 sky130_fd_sc_hd__dfrtn_1_27/a_1462_47# RESET_COUNTERn 0.00fF
C274 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_448_47# -0.00fF
C275 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# -0.00fF
C276 sky130_fd_sc_hd__o211a_1_0/a_79_21# out 0.01fF
C277 sky130_fd_sc_hd__o311a_1_0/a_266_47# SEL_CONV_TIME[2] 0.00fF
C278 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C279 sky130_fd_sc_hd__nor3_1_4/A sky130_fd_sc_hd__inv_1_6/A 0.01fF
C280 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C281 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C282 sky130_fd_sc_hd__mux4_2_0/a_788_316# SEL_CONV_TIME[2] 0.00fF
C283 sky130_fd_sc_hd__dfrtn_1_23/a_651_413# VDD 0.00fF
C284 sky130_fd_sc_hd__dfrtn_1_12/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C285 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C286 sky130_fd_sc_hd__dfrtn_1_30/a_805_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C287 sky130_fd_sc_hd__nor3_2_0/a_281_297# sky130_fd_sc_hd__dfrtn_1_12/a_639_47# 0.00fF
C288 DOUT[13] sky130_fd_sc_hd__dfrtn_1_30/a_1270_413# 0.00fF
C289 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_651_413# 0.00fF
C290 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C291 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C292 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C293 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_38/a_761_289# 0.00fF
C294 sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# DOUT[2] 0.00fF
C295 sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# sky130_fd_sc_hd__mux4_2_0/a_872_316# 0.00fF
C296 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C297 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__o311a_1_0/A3 0.01fF
C298 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_3/a_27_47# 0.00fF
C299 sky130_fd_sc_hd__dfrtn_1_7/a_543_47# VDD 0.03fF
C300 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# DOUT[14] 0.15fF
C301 sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# RESET_COUNTERn 0.02fF
C302 sky130_fd_sc_hd__dfrtn_1_36/a_639_47# DOUT[21] 0.00fF
C303 sky130_fd_sc_hd__dfrtn_1_37/a_639_47# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C304 sky130_fd_sc_hd__dfrtn_1_3/a_761_289# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C305 sky130_fd_sc_hd__inv_1_9/A RESET_COUNTERn 0.17fF
C306 DOUT[4] sky130_fd_sc_hd__dfrtn_1_28/a_761_289# 0.00fF
C307 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# sky130_fd_sc_hd__or2_2_0/B 0.01fF
C308 sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C309 sky130_fd_sc_hd__o311a_1_0/a_266_297# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C310 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C311 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C312 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# VDD 0.00fF
C313 VDD DOUT[20] 0.57fF
C314 sky130_fd_sc_hd__dfrtn_1_11/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C315 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C316 sky130_fd_sc_hd__dfrtn_1_18/a_193_47# sky130_fd_sc_hd__inv_1_35/A 0.01fF
C317 sky130_fd_sc_hd__nand2_1_2/a_113_47# RESET_COUNTERn 0.00fF
C318 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# -0.00fF
C319 sky130_fd_sc_hd__inv_1_15/A sky130_fd_sc_hd__inv_1_6/A 0.01fF
C320 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__dfrtn_1_25/a_639_47# 0.00fF
C321 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__inv_1_22/A 0.01fF
C322 sky130_fd_sc_hd__dfrtn_1_21/a_193_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C323 sky130_fd_sc_hd__dfrtn_1_18/a_1217_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C324 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C325 sky130_fd_sc_hd__nor3_1_7/a_193_297# RESET_COUNTERn 0.00fF
C326 sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# DOUT[23] 0.00fF
C327 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# 0.00fF
C328 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# 0.00fF
C329 sky130_fd_sc_hd__or3_1_0/a_111_297# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C330 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# 0.00fF
C331 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# SEL_CONV_TIME[1] 0.00fF
C332 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# 0.00fF
C333 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# 0.00fF
C334 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# sky130_fd_sc_hd__dfrtn_1_27/a_761_289# 0.00fF
C335 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C336 sky130_fd_sc_hd__o2111a_2_0/a_386_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C337 sky130_fd_sc_hd__dfrtn_1_26/a_543_47# sky130_fd_sc_hd__dfrtn_1_38/a_1462_47# 0.00fF
C338 CLK_REF sky130_fd_sc_hd__o211a_1_1/X 0.00fF
C339 sky130_fd_sc_hd__dfrtn_1_42/a_543_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C340 sky130_fd_sc_hd__dfrtn_1_27/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C341 sky130_fd_sc_hd__dfrtn_1_8/a_1217_47# VDD 0.00fF
C342 sky130_fd_sc_hd__dfrtn_1_8/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C343 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__inv_1_5/Y 0.02fF
C344 sky130_fd_sc_hd__dfrtn_1_34/a_448_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C345 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_805_47# -0.00fF
C346 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C347 DOUT[13] sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# 0.00fF
C348 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C349 sky130_fd_sc_hd__dfrtn_1_24/a_805_47# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C350 sky130_fd_sc_hd__dfrtn_1_32/a_27_47# RESET_COUNTERn 0.00fF
C351 sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# DOUT[21] 0.00fF
C352 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__dfrtn_1_34/a_761_289# 0.00fF
C353 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__dfrtn_1_34/a_543_47# 0.00fF
C354 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C355 sky130_fd_sc_hd__or3b_2_0/B SEL_CONV_TIME[1] 0.44fF
C356 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__inv_1_45/A 0.00fF
C357 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# CLK_REF 0.02fF
C358 sky130_fd_sc_hd__dfrtn_1_19/a_543_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C359 DOUT[4] sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# 0.00fF
C360 sky130_fd_sc_hd__dfrtn_1_31/a_1462_47# SEL_CONV_TIME[0] 0.00fF
C361 sky130_fd_sc_hd__o311a_1_0/a_368_297# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C362 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__dfrtn_1_22/a_193_47# -0.29fF
C363 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__inv_1_1/Y 0.00fF
C364 sky130_fd_sc_hd__dfrtn_1_36/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C365 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_15/a_27_47# 0.00fF
C366 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C367 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__or2b_1_0/X 0.17fF
C368 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C369 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C370 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C371 sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C372 sky130_fd_sc_hd__dfrtn_1_25/a_651_413# sky130_fd_sc_hd__or3_1_0/C 0.01fF
C373 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.04fF
C374 sky130_fd_sc_hd__nor3_2_0/a_27_297# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C375 sky130_fd_sc_hd__dfrtn_1_39/a_543_47# sky130_fd_sc_hd__inv_1_32/A 0.01fF
C376 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__mux4_2_0/a_872_316# 0.01fF
C377 sky130_fd_sc_hd__dfrtn_1_7/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C378 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# 0.00fF
C379 sky130_fd_sc_hd__dfrtn_1_17/a_1270_413# RESET_COUNTERn 0.00fF
C380 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# DOUT[14] 0.00fF
C381 sky130_fd_sc_hd__dfrtn_1_41/a_651_413# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C382 sky130_fd_sc_hd__dfrtn_1_9/a_805_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C383 DOUT[7] DOUT[14] 0.10fF
C384 sky130_fd_sc_hd__nor2_1_0/a_109_297# RESET_COUNTERn 0.00fF
C385 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__inv_1_7/A 0.01fF
C386 sky130_fd_sc_hd__dfrtn_1_19/a_27_47# sky130_fd_sc_hd__inv_1_34/Y 0.01fF
C387 sky130_fd_sc_hd__dfrtn_1_0/a_448_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C388 DOUT[4] sky130_fd_sc_hd__dfrtn_1_35/a_761_289# 0.01fF
C389 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C390 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C391 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_2/a_543_47# 0.00fF
C392 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_639_47# 0.00fF
C393 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# 0.00fF
C394 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C395 sky130_fd_sc_hd__dfrtn_1_31/a_448_47# RESET_COUNTERn 0.01fF
C396 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C397 sky130_fd_sc_hd__dfrtn_1_20/a_651_413# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C398 sky130_fd_sc_hd__inv_1_9/Y DOUT[21] 0.21fF
C399 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_12/a_193_47# 0.00fF
C400 sky130_fd_sc_hd__dfrtn_1_9/a_448_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C401 sky130_fd_sc_hd__or2_2_0/a_39_297# sky130_fd_sc_hd__dfrtn_1_19/a_448_47# 0.00fF
C402 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# SEL_CONV_TIME[1] 0.00fF
C403 sky130_fd_sc_hd__inv_1_2/A DOUT[3] 0.16fF
C404 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C405 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# 0.00fF
C406 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_8/a_27_47# 0.02fF
C407 sky130_fd_sc_hd__inv_1_31/Y sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C408 sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# DOUT[2] 0.01fF
C409 sky130_fd_sc_hd__inv_1_12/A DOUT[14] 0.01fF
C410 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# sky130_fd_sc_hd__dfrtn_1_23/a_193_47# 0.00fF
C411 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__dfrtn_1_23/a_761_289# 0.00fF
C412 sky130_fd_sc_hd__dfrtn_1_22/a_761_289# sky130_fd_sc_hd__dfrtn_1_23/a_27_47# 0.00fF
C413 sky130_fd_sc_hd__dfrtn_1_31/a_1283_21# DONE 0.00fF
C414 sky130_fd_sc_hd__mux4_2_0/a_872_316# sky130_fd_sc_hd__inv_1_33/A 0.01fF
C415 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_21/a_448_47# 0.01fF
C416 sky130_fd_sc_hd__dfrtn_1_9/a_543_47# sky130_fd_sc_hd__inv_1_37/A 0.01fF
C417 sky130_fd_sc_hd__dfrtn_1_38/a_193_47# sky130_fd_sc_hd__inv_1_27/Y 0.13fF
C418 sky130_fd_sc_hd__dfrtn_1_5/a_805_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C419 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C420 sky130_fd_sc_hd__dfrtn_1_29/a_639_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C421 sky130_fd_sc_hd__dfrtn_1_23/a_1462_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C422 sky130_fd_sc_hd__dfrtn_1_32/a_1217_47# RESET_COUNTERn 0.00fF
C423 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# SEL_CONV_TIME[0] 0.00fF
C424 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_33/a_651_413# 0.00fF
C425 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__dfrtn_1_33/a_761_289# 0.00fF
C426 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__dfrtn_1_33/a_543_47# 0.00fF
C427 sky130_fd_sc_hd__o311a_1_0/a_266_47# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C428 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# RESET_COUNTERn 0.01fF
C429 sky130_fd_sc_hd__dfrtn_1_8/a_805_47# sky130_fd_sc_hd__inv_1_9/Y 0.00fF
C430 sky130_fd_sc_hd__dfrtn_1_28/a_639_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C431 sky130_fd_sc_hd__inv_1_39/A sky130_fd_sc_hd__inv_1_39/Y 0.02fF
C432 sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C433 sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# outb 0.00fF
C434 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# 0.00fF
C435 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__o211a_1_1/X 0.00fF
C436 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# VDD 0.17fF
C437 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C438 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C439 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_3/A 0.02fF
C440 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C441 sky130_fd_sc_hd__dfrtn_1_37/a_805_47# VDD 0.00fF
C442 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__inv_1_14/A 0.10fF
C443 sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__inv_1_46/Y 0.00fF
C444 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# 0.00fF
C445 sky130_fd_sc_hd__inv_1_44/Y sky130_fd_sc_hd__inv_1_48/A 0.02fF
C446 sky130_fd_sc_hd__dfrtn_1_3/a_639_47# VDD 0.00fF
C447 sky130_fd_sc_hd__dfrtn_1_3/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C448 sky130_fd_sc_hd__dfrtn_1_14/a_651_413# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C449 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__inv_1_35/A 0.01fF
C450 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# 0.00fF
C451 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# 0.00fF
C452 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__dfrtp_1_2/a_761_289# 0.00fF
C453 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__dfrtp_1_2/a_543_47# 0.00fF
C454 sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C455 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C456 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C457 sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# RESET_COUNTERn 0.00fF
C458 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C459 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C460 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C461 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C462 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# 0.00fF
C463 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C464 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.01fF
C465 sky130_fd_sc_hd__nor3_1_2/a_109_297# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C466 sky130_fd_sc_hd__dfrtn_1_42/a_193_47# VDD 0.10fF
C467 DOUT[1] sky130_fd_sc_hd__inv_1_36/A 0.78fF
C468 sky130_fd_sc_hd__dfrtn_1_36/a_1270_413# sky130_fd_sc_hd__inv_1_38/A 0.00fF
C469 sky130_fd_sc_hd__dfrtn_1_19/a_1217_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C470 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# DOUT[21] 0.00fF
C471 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# RESET_COUNTERn 0.28fF
C472 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__inv_1_8/A 0.01fF
C473 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.01fF
C474 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__dfrtn_1_23/a_543_47# -0.00fF
C475 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C476 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__nor3_1_3/a_193_297# 0.00fF
C477 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C478 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C479 VDD sky130_fd_sc_hd__inv_1_38/A 0.54fF
C480 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# VDD 0.04fF
C481 sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C482 sky130_fd_sc_hd__dfrtn_1_4/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C483 sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# VDD 0.07fF
C484 sky130_fd_sc_hd__dfrtn_1_14/a_543_47# DOUT[11] 0.00fF
C485 sky130_fd_sc_hd__dfrtn_1_38/a_543_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C486 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_37/a_448_47# 0.00fF
C487 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C488 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# 0.00fF
C489 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# 0.00fF
C490 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# 0.01fF
C491 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.00fF
C492 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_26/a_651_413# 0.00fF
C493 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__dfrtn_1_26/a_805_47# 0.00fF
C494 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__dfrtn_1_26/a_639_47# 0.00fF
C495 sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C496 sky130_fd_sc_hd__dfrtn_1_7/a_543_47# DOUT[3] 0.00fF
C497 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_29/a_543_47# 0.00fF
C498 sky130_fd_sc_hd__dfrtn_1_25/a_1462_47# SEL_CONV_TIME[1] 0.00fF
C499 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C500 sky130_fd_sc_hd__dfrtn_1_21/a_193_47# VDD 0.08fF
C501 sky130_fd_sc_hd__inv_1_31/A SEL_CONV_TIME[1] 0.09fF
C502 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_8/a_1217_47# 0.00fF
C503 sky130_fd_sc_hd__dfrtn_1_19/a_1270_413# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C504 sky130_fd_sc_hd__o211a_1_1/a_510_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C505 sky130_fd_sc_hd__dfrtn_1_16/a_193_47# sky130_fd_sc_hd__dfrtn_1_16/a_651_413# -0.00fF
C506 sky130_fd_sc_hd__dfrtn_1_7/a_543_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C507 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# DOUT[3] 0.00fF
C508 DOUT[20] DOUT[3] 0.28fF
C509 sky130_fd_sc_hd__o311a_1_0/a_266_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C510 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# sky130_fd_sc_hd__o311a_1_0/A3 0.01fF
C511 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_193_47# 0.01fF
C512 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__dfrtn_1_7/a_27_47# 0.01fF
C513 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__nor3_1_4/A 0.01fF
C514 sky130_fd_sc_hd__inv_1_27/A RESET_COUNTERn 0.19fF
C515 sky130_fd_sc_hd__nor3_1_20/a_193_297# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C516 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__nor3_1_4/a_193_297# 0.00fF
C517 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__nor3_1_4/a_109_297# 0.00fF
C518 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_3/a_543_47# 0.00fF
C519 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# 0.05fF
C520 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C521 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__inv_1_38/Y 0.26fF
C522 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C523 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__inv_1_32/Y 0.01fF
C524 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__dfrtn_1_28/a_1108_47# -0.00fF
C525 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__dfrtn_1_16/a_651_413# 0.00fF
C526 sky130_fd_sc_hd__nor3_2_2/a_281_297# sky130_fd_sc_hd__dfrtn_1_16/a_448_47# 0.00fF
C527 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__dfrtn_1_33/a_639_47# 0.00fF
C528 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# VDD 0.05fF
C529 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C530 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C531 sky130_fd_sc_hd__inv_1_2/A DOUT[20] 0.57fF
C532 sky130_fd_sc_hd__dfrtp_1_1/a_639_47# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C533 sky130_fd_sc_hd__dfrtp_1_3/a_1217_47# RESET_COUNTERn 0.00fF
C534 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1_6/a_651_413# -0.00fF
C535 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__dfrtn_1_6/a_448_47# -0.00fF
C536 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__o211a_1_1/a_510_47# 0.00fF
C537 sky130_fd_sc_hd__dfrtp_1_1/a_805_47# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.00fF
C538 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C539 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C540 sky130_fd_sc_hd__dfrtn_1_22/a_761_289# RESET_COUNTERn 0.00fF
C541 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_448_47# 0.00fF
C542 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C543 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C544 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C545 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C546 sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# VDD 0.11fF
C547 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C548 sky130_fd_sc_hd__dfrtn_1_25/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C549 sky130_fd_sc_hd__dfrtn_1_25/a_1217_47# VDD 0.00fF
C550 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__dfrtn_1_3/a_27_47# 0.00fF
C551 sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# sky130_fd_sc_hd__dfrtn_1_3/a_761_289# 0.00fF
C552 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__dfrtn_1_3/a_543_47# 0.00fF
C553 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_3/a_651_413# 0.00fF
C554 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__dfrtn_1_3/a_193_47# 0.00fF
C555 sky130_fd_sc_hd__dfrtn_1_41/a_1270_413# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C556 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_805_47# 0.00fF
C557 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# 0.00fF
C558 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_3/a_639_47# 0.00fF
C559 sky130_fd_sc_hd__nor3_1_11/a_109_297# VIN 0.00fF
C560 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C561 sky130_fd_sc_hd__o221ai_1_0/a_109_47# SEL_CONV_TIME[1] 0.00fF
C562 VDD sky130_fd_sc_hd__inv_1_11/Y 0.62fF
C563 sky130_fd_sc_hd__nor3_2_3/a_27_297# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C564 sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# VDD 0.13fF
C565 sky130_fd_sc_hd__dfrtn_1_20/a_805_47# sky130_fd_sc_hd__inv_1_35/Y 0.00fF
C566 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__dfrtn_1_25/a_543_47# 0.00fF
C567 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__o221ai_1_0/a_295_297# 0.00fF
C568 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__inv_1_5/Y 0.01fF
C569 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_5/A 0.00fF
C570 sky130_fd_sc_hd__inv_1_33/A SEL_CONV_TIME[1] 0.06fF
C571 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_40/Y 0.02fF
C572 sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# sky130_fd_sc_hd__inv_1_1/A 0.01fF
C573 sky130_fd_sc_hd__dfrtn_1_41/a_448_47# DOUT[2] 0.00fF
C574 sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# 0.00fF
C575 sky130_fd_sc_hd__dfrtp_1_1/a_639_47# sky130_fd_sc_hd__dfrtp_1_2/a_651_413# 0.00fF
C576 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# 0.00fF
C577 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C578 sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C579 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C580 sky130_fd_sc_hd__dfrtn_1_17/a_193_47# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C581 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C582 sky130_fd_sc_hd__dfrtn_1_42/a_1462_47# VDD 0.00fF
C583 sky130_fd_sc_hd__dfrtn_1_42/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C584 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# 0.00fF
C585 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# RESET_COUNTERn 0.02fF
C586 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# DOUT[14] 0.00fF
C587 sky130_fd_sc_hd__dfrtn_1_17/a_193_47# sky130_fd_sc_hd__inv_1_29/Y 0.00fF
C588 sky130_fd_sc_hd__dfrtn_1_8/a_193_47# DOUT[21] 0.02fF
C589 VDD sky130_fd_sc_hd__inv_1_3/Y 0.43fF
C590 sky130_fd_sc_hd__nor3_1_6/a_109_297# RESET_COUNTERn 0.00fF
C591 VDD sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.07fF
C592 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_20/a_193_47# -0.33fF
C593 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C594 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C595 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C596 sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# RESET_COUNTERn 0.00fF
C597 sky130_fd_sc_hd__nand3b_1_1/Y RESET_COUNTERn 0.01fF
C598 sky130_fd_sc_hd__dfrtn_1_38/a_543_47# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C599 sky130_fd_sc_hd__dfrtn_1_10/a_1217_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C600 sky130_fd_sc_hd__dfrtn_1_41/a_1270_413# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C601 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__dfrtn_1_38/a_543_47# 0.00fF
C602 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C603 sky130_fd_sc_hd__dfrtn_1_41/a_651_413# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C604 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_651_413# 0.00fF
C605 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_36/a_1462_47# 0.00fF
C606 sky130_fd_sc_hd__dfrtn_1_19/a_27_47# VDD 0.18fF
C607 sky130_fd_sc_hd__dfrtp_1_3/a_543_47# DOUT[23] 0.00fF
C608 DOUT[9] sky130_fd_sc_hd__nor3_1_4/a_109_297# 0.00fF
C609 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C610 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__or2b_1_0/a_219_297# 0.00fF
C611 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_1/a_543_47# 0.00fF
C612 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_1/a_448_47# 0.00fF
C613 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_1/a_27_47# 0.00fF
C614 VDD sky130_fd_sc_hd__inv_1_29/Y 0.09fF
C615 sky130_fd_sc_hd__o311a_1_0/a_585_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C616 sky130_fd_sc_hd__o221ai_1_0/a_493_297# VDD 0.00fF
C617 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__mux4_2_0/a_872_316# 0.01fF
C618 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.08fF
C619 sky130_fd_sc_hd__mux4_2_0/a_600_345# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C620 sky130_fd_sc_hd__inv_1_50/A SEL_CONV_TIME[0] 0.15fF
C621 sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C622 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# SEL_CONV_TIME[1] 0.01fF
C623 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_448_47# -0.00fF
C624 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# -0.00fF
C625 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__o221ai_1_0/a_295_297# 0.00fF
C626 sky130_fd_sc_hd__dfrtp_1_3/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C627 sky130_fd_sc_hd__dfrtn_1_33/a_651_413# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C628 sky130_fd_sc_hd__dfrtn_1_16/a_1270_413# DOUT[15] 0.00fF
C629 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C630 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C631 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__inv_1_5/Y 0.01fF
C632 sky130_fd_sc_hd__dfrtn_1_23/a_1270_413# DOUT[21] 0.00fF
C633 sky130_fd_sc_hd__dfrtn_1_23/a_543_47# RESET_COUNTERn 0.01fF
C634 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C635 sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C636 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__dfrtn_1_26/a_448_47# 0.00fF
C637 sky130_fd_sc_hd__nor3_1_0/A RESET_COUNTERn 0.02fF
C638 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# sky130_fd_sc_hd__dfrtn_1_7/a_805_47# 0.00fF
C639 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__dfrtn_1_7/a_1217_47# 0.00fF
C640 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_1462_47# 0.00fF
C641 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# sky130_fd_sc_hd__dfrtn_1_7/a_27_47# 0.00fF
C642 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# 0.00fF
C643 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__dfrtn_1_7/a_651_413# 0.00fF
C644 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# sky130_fd_sc_hd__dfrtn_1_7/a_761_289# 0.00fF
C645 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# sky130_fd_sc_hd__dfrtn_1_7/a_193_47# 0.00fF
C646 sky130_fd_sc_hd__dfrtn_1_12/a_1270_413# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C647 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# DOUT[6] 0.00fF
C648 sky130_fd_sc_hd__dfrtn_1_7/a_543_47# DOUT[20] 0.01fF
C649 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# DOUT[7] 0.02fF
C650 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# DOUT[8] 0.00fF
C651 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C652 sky130_fd_sc_hd__dfrtp_1_0/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C653 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# sky130_fd_sc_hd__dfrtn_1_0/a_1462_47# 0.00fF
C654 sky130_fd_sc_hd__inv_1_51/Y RESET_COUNTERn 0.01fF
C655 sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# 0.00fF
C656 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_0/a_761_289# -0.00fF
C657 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# DOUT[7] 0.00fF
C658 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# RESET_COUNTERn 0.00fF
C659 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# DOUT[6] 0.00fF
C660 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# DOUT[20] 0.00fF
C661 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C662 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C663 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_5/a_805_47# 0.00fF
C664 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# 0.00fF
C665 sky130_fd_sc_hd__inv_1_36/Y sky130_fd_sc_hd__nor3_2_3/C 0.08fF
C666 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# SEL_CONV_TIME[2] 0.00fF
C667 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__mux4_1_0/a_247_21# -0.00fF
C668 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__mux4_1_0/a_277_47# -0.00fF
C669 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_32/a_1270_413# 0.00fF
C670 CLK_REF sky130_fd_sc_hd__dfrtn_1_20/a_805_47# 0.00fF
C671 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C672 sky130_fd_sc_hd__dfrtn_1_27/a_193_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C673 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_543_47# 0.00fF
C674 sky130_fd_sc_hd__dfrtn_1_26/a_761_289# sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.00fF
C675 sky130_fd_sc_hd__dfrtn_1_26/a_543_47# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C676 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# 0.00fF
C677 sky130_fd_sc_hd__dfrtn_1_30/a_805_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C678 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C679 sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# VDD 0.11fF
C680 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_10/a_1217_47# -0.00fF
C681 sky130_fd_sc_hd__o2111a_2_0/a_386_47# sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.00fF
C682 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__inv_1_32/A 0.01fF
C683 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__o311a_1_0/a_368_297# 0.00fF
C684 sky130_fd_sc_hd__inv_1_49/Y VDD 0.38fF
C685 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# outb 0.00fF
C686 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# SEL_CONV_TIME[0] 0.00fF
C687 sky130_fd_sc_hd__dfrtn_1_29/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C688 sky130_fd_sc_hd__inv_1_34/Y sky130_fd_sc_hd__inv_1_28/A 0.03fF
C689 sky130_fd_sc_hd__inv_1_54/Y RESET_COUNTERn 0.12fF
C690 en DOUT[14] 0.03fF
C691 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__dfrtn_1_3/a_193_47# 0.00fF
C692 sky130_fd_sc_hd__nor3_1_3/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C693 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__or2_2_0/B 0.00fF
C694 sky130_fd_sc_hd__dfrtn_1_9/a_543_47# DOUT[14] 0.00fF
C695 sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C696 sky130_fd_sc_hd__dfrtn_1_17/a_1462_47# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C697 sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# sky130_fd_sc_hd__dfrtn_1_19/a_651_413# 0.00fF
C698 DOUT[15] RESET_COUNTERn 0.05fF
C699 sky130_fd_sc_hd__dfrtn_1_26/a_651_413# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C700 sky130_fd_sc_hd__dfrtn_1_16/a_1217_47# RESET_COUNTERn 0.00fF
C701 sky130_fd_sc_hd__dfrtn_1_8/a_1462_47# DOUT[21] 0.00fF
C702 sky130_fd_sc_hd__dfrtn_1_8/a_651_413# RESET_COUNTERn 0.00fF
C703 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__inv_1_38/A 0.01fF
C704 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# sky130_fd_sc_hd__o211a_1_0/X 0.00fF
C705 sky130_fd_sc_hd__dfrtn_1_9/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C706 sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# SEL_CONV_TIME[1] 0.05fF
C707 VDD sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# 0.00fF
C708 sky130_fd_sc_hd__inv_1_27/A SEL_CONV_TIME[2] 0.00fF
C709 sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C710 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C711 sky130_fd_sc_hd__dfrtn_1_32/a_448_47# sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C712 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# 0.01fF
C713 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_30/a_193_47# 0.01fF
C714 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_30/a_761_289# 0.00fF
C715 sky130_fd_sc_hd__dfrtn_1_19/a_1217_47# VDD 0.00fF
C716 sky130_fd_sc_hd__nor3_1_8/a_193_297# VDD 0.00fF
C717 sky130_fd_sc_hd__nor3_2_3/B DOUT[18] 0.14fF
C718 sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C719 sky130_fd_sc_hd__inv_1_21/Y DOUT[12] 0.00fF
C720 sky130_fd_sc_hd__dfrtn_1_11/a_761_289# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C721 sky130_fd_sc_hd__or2b_1_0/a_301_297# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C722 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C723 sky130_fd_sc_hd__dfrtn_1_31/a_639_47# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C724 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_27/a_1270_413# 0.00fF
C725 sky130_fd_sc_hd__nand3b_1_1/Y SEL_CONV_TIME[3] 0.02fF
C726 DOUT[4] sky130_fd_sc_hd__dfrtn_1_36/a_1270_413# 0.00fF
C727 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C728 sky130_fd_sc_hd__nor3_1_10/a_109_297# sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# 0.00fF
C729 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# 0.00fF
C730 sky130_fd_sc_hd__dfrtn_1_34/a_448_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C731 sky130_fd_sc_hd__dfrtn_1_22/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C732 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C733 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__inv_1_47/Y 0.00fF
C734 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# 0.00fF
C735 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_1/Y 0.00fF
C736 VDD sky130_fd_sc_hd__inv_1_0/Y 0.51fF
C737 sky130_fd_sc_hd__dfrtn_1_7/a_1462_47# DOUT[7] 0.00fF
C738 sky130_fd_sc_hd__dfrtn_1_7/a_805_47# RESET_COUNTERn 0.00fF
C739 DOUT[4] VDD 5.28fF
C740 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C741 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# DOUT[3] 0.00fF
C742 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__nand2_1_1/a_113_47# 0.00fF
C743 sky130_fd_sc_hd__dfrtn_1_30/a_543_47# VDD 0.07fF
C744 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C745 sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# DOUT[3] 0.00fF
C746 SEL_CONV_TIME[1] sky130_fd_sc_hd__o2111a_2_0/X 0.03fF
C747 sky130_fd_sc_hd__inv_1_15/A sky130_fd_sc_hd__inv_1_8/A 0.00fF
C748 sky130_fd_sc_hd__dfrtn_1_16/a_543_47# DOUT[23] 0.00fF
C749 sky130_fd_sc_hd__or3b_2_0/B DOUT[21] 0.00fF
C750 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__inv_1_48/A 0.01fF
C751 sky130_fd_sc_hd__dfrtn_1_30/a_761_289# sky130_fd_sc_hd__dfrtn_1_31/a_27_47# 0.01fF
C752 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__dfrtn_1_31/a_193_47# 0.00fF
C753 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_761_289# 0.01fF
C754 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# DOUT[14] 0.01fF
C755 sky130_fd_sc_hd__nor3_1_1/a_109_297# RESET_COUNTERn 0.00fF
C756 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# sky130_fd_sc_hd__inv_1_15/A 0.01fF
C757 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__dfrtn_1_35/a_1108_47# -0.00fF
C758 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__inv_1_2/A 0.01fF
C759 sky130_fd_sc_hd__dfrtp_1_1/a_639_47# CLK_REF 0.00fF
C760 sky130_fd_sc_hd__mux4_2_0/X SEL_CONV_TIME[1] 0.08fF
C761 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C762 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C763 sky130_fd_sc_hd__nor3_1_3/a_193_297# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C764 sky130_fd_sc_hd__dfrtn_1_20/a_1270_413# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C765 sky130_fd_sc_hd__dfrtn_1_14/a_651_413# DOUT[17] 0.00fF
C766 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_1478_413# -0.00fF
C767 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_668_97# -0.00fF
C768 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__inv_1_11/Y 0.01fF
C769 sky130_fd_sc_hd__nand3b_1_1/Y SEL_CONV_TIME[2] 0.00fF
C770 sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# sky130_fd_sc_hd__dfrtn_1_27/a_448_47# 0.00fF
C771 sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# sky130_fd_sc_hd__dfrtn_1_27/a_543_47# 0.00fF
C772 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# sky130_fd_sc_hd__dfrtn_1_27/a_805_47# 0.00fF
C773 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C774 sky130_fd_sc_hd__o211a_1_1/a_297_297# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C775 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# SEL_CONV_TIME[1] 0.01fF
C776 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C777 sky130_fd_sc_hd__dfrtn_1_40/a_1462_47# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C778 sky130_fd_sc_hd__dfrtn_1_16/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C779 sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C780 sky130_fd_sc_hd__dfrtn_1_5/a_805_47# VDD 0.00fF
C781 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# SEL_CONV_TIME[0] 0.00fF
C782 sky130_fd_sc_hd__dfrtn_1_8/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C783 sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C784 sky130_fd_sc_hd__dfrtn_1_37/a_1462_47# SEL_CONV_TIME[0] 0.00fF
C785 sky130_fd_sc_hd__nand3b_1_0/a_232_47# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C786 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# sky130_fd_sc_hd__dfrtn_1_11/a_27_47# 0.00fF
C787 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_761_289# 0.00fF
C788 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_11/a_193_47# 0.00fF
C789 sky130_fd_sc_hd__o211a_1_1/a_79_21# VDD 0.08fF
C790 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C791 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_12/a_448_47# 0.00fF
C792 DOUT[4] sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# 0.00fF
C793 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C794 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__o211a_1_1/X 0.01fF
C795 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__nor3_1_5/A 0.00fF
C796 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__o311a_1_0/A3 0.01fF
C797 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C798 sky130_fd_sc_hd__inv_1_47/Y VDD 0.28fF
C799 sky130_fd_sc_hd__dfrtn_1_33/a_805_47# SEL_CONV_TIME[1] 0.00fF
C800 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__dfrtn_1_40/a_761_289# 0.00fF
C801 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__dfrtn_1_40/a_193_47# 0.00fF
C802 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_17/a_761_289# 0.00fF
C803 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_651_413# 0.00fF
C804 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_448_47# 0.00fF
C805 sky130_fd_sc_hd__dfrtp_1_2/a_448_47# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C806 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C807 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# 0.00fF
C808 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__dfrtn_1_14/a_193_47# 0.00fF
C809 sky130_fd_sc_hd__dfrtn_1_12/a_761_289# sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# 0.00fF
C810 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_14/a_651_413# 0.00fF
C811 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C812 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_14/a_193_47# 0.02fF
C813 sky130_fd_sc_hd__nor3_2_2/a_281_297# sky130_fd_sc_hd__dfrtn_1_42/a_543_47# 0.00fF
C814 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C815 sky130_fd_sc_hd__dfrtn_1_23/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C816 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# sky130_fd_sc_hd__inv_1_6/A 0.01fF
C817 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# DOUT[14] 0.01fF
C818 sky130_fd_sc_hd__nor3_1_13/a_193_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C819 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# 0.00fF
C820 sky130_fd_sc_hd__dfrtp_1_2/a_448_47# VDD 0.01fF
C821 DOUT[19] sky130_fd_sc_hd__inv_1_3/A 0.03fF
C822 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C823 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C824 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# sky130_fd_sc_hd__o221ai_1_0/a_493_297# 0.00fF
C825 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C826 sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C827 DOUT[23] DOUT[21] 0.01fF
C828 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C829 sky130_fd_sc_hd__dfrtn_1_16/a_761_289# sky130_fd_sc_hd__inv_1_26/A 0.00fF
C830 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C831 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# VDD 0.00fF
C832 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# DOUT[21] 0.00fF
C833 sky130_fd_sc_hd__dfrtn_1_42/a_1270_413# sky130_fd_sc_hd__dfrtn_1_23/a_27_47# 0.00fF
C834 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C835 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_6/a_761_289# 0.00fF
C836 sky130_fd_sc_hd__dfrtn_1_38/a_1270_413# SEL_CONV_TIME[1] 0.00fF
C837 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C838 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__inv_1_1/A 0.02fF
C839 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# RESET_COUNTERn 0.01fF
C840 sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# sky130_fd_sc_hd__inv_1_48/Y 0.01fF
C841 sky130_fd_sc_hd__dfrtn_1_32/a_193_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C842 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C843 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C844 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C845 sky130_fd_sc_hd__dfrtn_1_11/a_1217_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C846 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__dfrtn_1_30/a_651_413# 0.00fF
C847 sky130_fd_sc_hd__inv_1_3/Y DOUT[3] 0.03fF
C848 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# DOUT[3] 0.00fF
C849 sky130_fd_sc_hd__dfrtn_1_33/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C850 sky130_fd_sc_hd__dfrtn_1_33/a_639_47# VDD -0.00fF
C851 sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# RESET_COUNTERn 0.02fF
C852 sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C853 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C854 VDD outb 5.14fF
C855 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_3/Y 0.02fF
C856 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C857 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# VDD 0.06fF
C858 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C859 sky130_fd_sc_hd__dfrtn_1_20/a_639_47# sky130_fd_sc_hd__inv_1_35/A 0.00fF
C860 sky130_fd_sc_hd__nor3_2_3/C DOUT[19] 0.18fF
C861 DOUT[22] sky130_fd_sc_hd__nor3_2_3/B 0.04fF
C862 sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C863 sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C864 sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# sky130_fd_sc_hd__inv_1_11/A 0.02fF
C865 sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# DOUT[14] 0.00fF
C866 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C867 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# sky130_fd_sc_hd__inv_1_15/A 0.01fF
C868 sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# DOUT[22] 0.00fF
C869 sky130_fd_sc_hd__inv_1_32/Y RESET_COUNTERn 0.04fF
C870 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# 0.00fF
C871 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# HEADER_0/a_508_138# 0.00fF
C872 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__or2_2_0/B 0.01fF
C873 DOUT[13] sky130_fd_sc_hd__dfrtn_1_36/a_543_47# 0.00fF
C874 sky130_fd_sc_hd__o211a_1_1/a_215_47# sky130_fd_sc_hd__dfrtn_1_17/a_805_47# 0.00fF
C875 sky130_fd_sc_hd__dfrtn_1_34/a_1217_47# SEL_CONV_TIME[1] 0.00fF
C876 sky130_fd_sc_hd__dfrtn_1_24/a_1270_413# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C877 sky130_fd_sc_hd__dfrtn_1_24/a_651_413# sky130_fd_sc_hd__dfrtn_1_29/a_761_289# 0.00fF
C878 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C879 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# sky130_fd_sc_hd__dfrtn_1_29/a_651_413# 0.00fF
C880 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_639_47# 0.00fF
C881 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# sky130_fd_sc_hd__dfrtn_1_29/a_448_47# 0.00fF
C882 sky130_fd_sc_hd__dfrtn_1_24/a_448_47# sky130_fd_sc_hd__dfrtn_1_29/a_543_47# 0.00fF
C883 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# 0.00fF
C884 sky130_fd_sc_hd__dfrtn_1_17/a_193_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C885 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# DOUT[6] 0.00fF
C886 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# DOUT[7] 0.01fF
C887 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# DOUT[20] 0.00fF
C888 sky130_fd_sc_hd__dfrtn_1_8/a_27_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C889 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# RESET_COUNTERn 0.32fF
C890 sky130_fd_sc_hd__nand3b_1_1/a_232_47# RESET_COUNTERn 0.00fF
C891 sky130_fd_sc_hd__or3_1_0/a_111_297# RESET_COUNTERn 0.00fF
C892 sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C893 sky130_fd_sc_hd__dfrtn_1_38/a_651_413# VDD 0.01fF
C894 sky130_fd_sc_hd__dfrtn_1_33/a_1108_47# sky130_fd_sc_hd__inv_1_45/A 0.00fF
C895 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# sky130_fd_sc_hd__dfrtn_1_11/a_1217_47# 0.00fF
C896 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__dfrtn_1_11/a_651_413# 0.00fF
C897 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__dfrtn_1_11/a_805_47# 0.00fF
C898 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_11/a_1462_47# 0.00fF
C899 sky130_fd_sc_hd__dfrtn_1_10/a_639_47# sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# 0.00fF
C900 sky130_fd_sc_hd__nor3_2_3/a_281_297# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C901 VDD sky130_fd_sc_hd__inv_1_28/A 0.48fF
C902 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C903 sky130_fd_sc_hd__dfrtn_1_42/a_1108_47# DOUT[15] 0.00fF
C904 sky130_fd_sc_hd__nor3_1_4/a_193_297# DOUT[19] 0.00fF
C905 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# 0.00fF
C906 sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# 0.00fF
C907 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/a_639_47# -0.00fF
C908 VIN DOUT[14] 1.35fF
C909 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_1/D 0.00fF
C910 sky130_fd_sc_hd__dfrtn_1_7/a_639_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C911 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# 0.00fF
C912 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__dfrtn_1_34/a_543_47# 0.00fF
C913 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_37/a_639_47# -0.00fF
C914 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__dfrtn_1_0/a_27_47# 0.01fF
C915 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# 0.01fF
C916 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C917 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# 0.00fF
C918 sky130_fd_sc_hd__nand2_1_2/Y RESET_COUNTERn 0.05fF
C919 sky130_fd_sc_hd__dfrtn_1_28/a_805_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C920 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C921 sky130_fd_sc_hd__dfrtn_1_26/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C922 sky130_fd_sc_hd__dfrtn_1_26/a_639_47# VDD 0.00fF
C923 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# DOUT[14] 0.00fF
C924 sky130_fd_sc_hd__nor3_1_10/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C925 sky130_fd_sc_hd__dfrtn_1_34/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C926 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__dfrtn_1_41/a_761_289# -0.00fF
C927 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_41/a_543_47# -0.00fF
C928 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C929 sky130_fd_sc_hd__dfrtn_1_34/a_805_47# VDD 0.00fF
C930 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_7/a_651_413# 0.00fF
C931 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C932 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_8/a_1283_21# 0.01fF
C933 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__inv_1_2/Y 0.10fF
C934 SLC_0/a_264_22# DOUT[15] 0.01fF
C935 sky130_fd_sc_hd__dfrtn_1_23/a_639_47# sky130_fd_sc_hd__inv_1_40/Y 0.00fF
C936 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_651_413# -0.00fF
C937 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_3/a_448_47# -0.00fF
C938 sky130_fd_sc_hd__o221ai_1_0/a_213_123# SEL_CONV_TIME[0] 0.01fF
C939 sky130_fd_sc_hd__inv_1_48/A sky130_fd_sc_hd__inv_1_48/Y 0.03fF
C940 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# RESET_COUNTERn 0.00fF
C941 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__inv_1_41/Y 0.07fF
C942 sky130_fd_sc_hd__dfrtn_1_25/a_651_413# RESET_COUNTERn 0.00fF
C943 sky130_fd_sc_hd__dfrtn_1_25/a_1462_47# DOUT[21] 0.00fF
C944 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__or2_2_0/a_121_297# 0.00fF
C945 sky130_fd_sc_hd__dfrtp_1_3/a_543_47# sky130_fd_sc_hd__or2_2_0/X 0.01fF
C946 sky130_fd_sc_hd__inv_1_4/A RESET_COUNTERn 0.17fF
C947 sky130_fd_sc_hd__dfrtn_1_32/a_1462_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C948 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C949 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# sky130_fd_sc_hd__inv_1_32/Y 0.00fF
C950 sky130_fd_sc_hd__inv_1_10/A DOUT[4] 0.00fF
C951 sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C952 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__o211a_1_1/a_510_47# 0.00fF
C953 sky130_fd_sc_hd__inv_1_25/A sky130_fd_sc_hd__nor3_2_3/C 0.03fF
C954 sky130_fd_sc_hd__dfrtn_1_18/a_27_47# RESET_COUNTERn 0.03fF
C955 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__inv_1_11/A 0.02fF
C956 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# DOUT[15] 0.00fF
C957 DOUT[15] DOUT[10] 0.03fF
C958 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# 0.01fF
C959 DOUT[4] sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# 0.00fF
C960 sky130_fd_sc_hd__nor3_1_8/a_193_297# DOUT[3] 0.00fF
C961 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C962 sky130_fd_sc_hd__nand3b_1_1/Y sky130_fd_sc_hd__or3_1_0/X 0.00fF
C963 sky130_fd_sc_hd__dfrtn_1_7/a_805_47# HEADER_0/a_508_138# 0.00fF
C964 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_543_47# 0.00fF
C965 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_761_289# 0.00fF
C966 sky130_fd_sc_hd__dfrtn_1_28/a_1283_21# SEL_CONV_TIME[1] 0.00fF
C967 sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C968 sky130_fd_sc_hd__dfrtn_1_42/a_1270_413# RESET_COUNTERn 0.00fF
C969 sky130_fd_sc_hd__mux4_2_0/a_1060_369# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C970 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__o311a_1_0/a_266_297# 0.00fF
C971 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C972 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C973 sky130_fd_sc_hd__inv_1_3/Y DOUT[20] 0.00fF
C974 DOUT[23] sky130_fd_sc_hd__dfrtp_1_1/D 0.09fF
C975 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_10/a_1270_413# 0.00fF
C976 sky130_fd_sc_hd__dfrtn_1_0/a_1462_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C977 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_639_47# 0.00fF
C978 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# sky130_fd_sc_hd__dfrtp_1_3/a_761_289# 0.00fF
C979 sky130_fd_sc_hd__dfrtp_1_2/a_639_47# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C980 sky130_fd_sc_hd__dfrtp_1_2/a_805_47# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C981 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C982 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C983 sky130_fd_sc_hd__nor3_1_2/a_193_297# DOUT[18] 0.00fF
C984 sky130_fd_sc_hd__dfrtn_1_17/a_1462_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C985 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C986 CLK_REF sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C987 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# RESET_COUNTERn 0.00fF
C988 sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# RESET_COUNTERn 0.00fF
C989 sky130_fd_sc_hd__dfrtn_1_24/a_448_47# SEL_CONV_TIME[0] 0.00fF
C990 sky130_fd_sc_hd__inv_1_37/A sky130_fd_sc_hd__inv_1_39/A 0.14fF
C991 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__inv_1_53/A 0.08fF
C992 VDD sky130_fd_sc_hd__nor3_2_3/A 0.67fF
C993 sky130_fd_sc_hd__inv_1_52/A RESET_COUNTERn 0.23fF
C994 sky130_fd_sc_hd__nor3_1_14/a_109_297# RESET_COUNTERn 0.00fF
C995 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__dfrtn_1_34/a_448_47# 0.00fF
C996 sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# RESET_COUNTERn 0.02fF
C997 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__inv_1_6/A 0.11fF
C998 sky130_fd_sc_hd__nor3_1_10/a_193_297# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C999 sky130_fd_sc_hd__inv_1_33/A DOUT[21] 0.00fF
C1000 sky130_fd_sc_hd__dfrtn_1_31/a_651_413# sky130_fd_sc_hd__inv_1_49/A 0.01fF
C1001 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C1002 DOUT[13] sky130_fd_sc_hd__dfrtn_1_31/a_1108_47# 0.00fF
C1003 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_761_289# 0.00fF
C1004 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_543_47# 0.01fF
C1005 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# SEL_CONV_TIME[2] 0.00fF
C1006 SLC_0/a_919_243# lc_out 0.00fF
C1007 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# 0.00fF
C1008 sky130_fd_sc_hd__dfrtn_1_28/a_543_47# VDD 0.06fF
C1009 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C1010 sky130_fd_sc_hd__nand3b_1_1/a_232_47# SEL_CONV_TIME[3] 0.00fF
C1011 sky130_fd_sc_hd__or3_1_0/a_111_297# SEL_CONV_TIME[3] 0.00fF
C1012 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# -0.00fF
C1013 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# sky130_fd_sc_hd__inv_1_7/Y 0.06fF
C1014 sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1015 sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C1016 sky130_fd_sc_hd__inv_1_0/Y DOUT[5] 0.00fF
C1017 sky130_fd_sc_hd__dfrtn_1_14/a_805_47# VDD 0.00fF
C1018 sky130_fd_sc_hd__dfrtn_1_12/a_1217_47# sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# 0.00fF
C1019 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__dfrtn_1_0/a_1217_47# 0.00fF
C1020 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_21/a_1217_47# 0.00fF
C1021 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C1022 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C1023 sky130_fd_sc_hd__dfrtp_1_0/a_805_47# RESET_COUNTERn 0.00fF
C1024 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C1025 sky130_fd_sc_hd__mux4_1_0/a_277_47# SEL_CONV_TIME[1] 0.06fF
C1026 sky130_fd_sc_hd__o221ai_1_0/a_109_47# sky130_fd_sc_hd__o311a_1_0/A3 0.01fF
C1027 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C1028 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# 0.00fF
C1029 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.02fF
C1030 sky130_fd_sc_hd__inv_1_1/A DOUT[14] 0.00fF
C1031 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C1032 lc_out out 0.19fF
C1033 sky130_fd_sc_hd__inv_1_2/Y DOUT[8] 0.00fF
C1034 sky130_fd_sc_hd__dfrtn_1_5/a_805_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C1035 sky130_fd_sc_hd__dfrtn_1_39/a_1217_47# RESET_COUNTERn 0.00fF
C1036 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C1037 sky130_fd_sc_hd__dfrtn_1_22/a_639_47# sky130_fd_sc_hd__inv_1_39/Y 0.00fF
C1038 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# VDD 0.09fF
C1039 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C1040 sky130_fd_sc_hd__inv_1_32/Y SEL_CONV_TIME[2] 0.01fF
C1041 sky130_fd_sc_hd__inv_1_33/A sky130_fd_sc_hd__o311a_1_0/A3 0.02fF
C1042 sky130_fd_sc_hd__dfrtn_1_42/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C1043 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# DOUT[21] 0.01fF
C1044 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# RESET_COUNTERn 0.01fF
C1045 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# sky130_fd_sc_hd__inv_1_42/A 0.01fF
C1046 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__o2111a_2_0/a_674_297# 0.00fF
C1047 sky130_fd_sc_hd__dfrtn_1_18/a_1217_47# RESET_COUNTERn 0.00fF
C1048 sky130_fd_sc_hd__inv_1_10/A outb 0.02fF
C1049 sky130_fd_sc_hd__dfrtp_1_3/a_1283_21# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C1050 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# 0.00fF
C1051 sky130_fd_sc_hd__or3b_2_0/X SEL_CONV_TIME[0] 0.11fF
C1052 sky130_fd_sc_hd__nand3b_1_1/Y sky130_fd_sc_hd__inv_1_53/A 0.00fF
C1053 DOUT[1] DOUT[16] 0.00fF
C1054 DOUT[1] sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C1055 DOUT[4] sky130_fd_sc_hd__dfrtn_1_8/a_27_47# 0.00fF
C1056 sky130_fd_sc_hd__inv_1_17/A sky130_fd_sc_hd__inv_1_22/A 0.00fF
C1057 sky130_fd_sc_hd__inv_1_24/A sky130_fd_sc_hd__inv_1_22/Y 0.00fF
C1058 VDD sky130_fd_sc_hd__inv_1_13/Y 0.30fF
C1059 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# SEL_CONV_TIME[0] 0.00fF
C1060 sky130_fd_sc_hd__dfrtn_1_23/a_543_47# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C1061 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1062 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_26/a_761_289# 0.00fF
C1063 sky130_fd_sc_hd__dfrtn_1_22/a_543_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C1064 sky130_fd_sc_hd__dfrtn_1_4/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1065 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# sky130_fd_sc_hd__dfrtn_1_42/a_761_289# -0.00fF
C1066 sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# SEL_CONV_TIME[0] 0.03fF
C1067 sky130_fd_sc_hd__dfrtn_1_3/a_639_47# sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C1068 sky130_fd_sc_hd__dfrtn_1_3/a_805_47# sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C1069 DOUT[13] sky130_fd_sc_hd__inv_1_52/Y 0.01fF
C1070 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1071 sky130_fd_sc_hd__mux4_1_0/a_247_21# VDD 0.04fF
C1072 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_7/Y 0.03fF
C1073 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# DOUT[3] 0.00fF
C1074 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C1075 SLC_0/a_919_243# sky130_fd_sc_hd__nor3_2_3/B 0.07fF
C1076 sky130_fd_sc_hd__dfrtn_1_10/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C1077 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# VDD 0.01fF
C1078 sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# RESET_COUNTERn 0.00fF
C1079 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# sky130_fd_sc_hd__dfrtn_1_15/a_193_47# 0.00fF
C1080 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C1081 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_543_47# 0.00fF
C1082 sky130_fd_sc_hd__dfrtp_1_0/a_761_289# DOUT[23] 0.00fF
C1083 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C1084 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C1085 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__o221ai_1_0/a_295_297# 0.00fF
C1086 sky130_fd_sc_hd__dfrtn_1_19/a_651_413# RESET_COUNTERn 0.01fF
C1087 sky130_fd_sc_hd__nor3_1_8/a_193_297# DOUT[20] 0.00fF
C1088 sky130_fd_sc_hd__nor3_1_8/a_109_297# DOUT[6] -0.00fF
C1089 sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C1090 CLK_REF sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# 0.00fF
C1091 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C1092 sky130_fd_sc_hd__mux4_2_0/a_1060_369# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C1093 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C1094 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_543_47# -0.00fF
C1095 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# -0.00fF
C1096 sky130_fd_sc_hd__mux4_2_0/a_372_413# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C1097 sky130_fd_sc_hd__dfrtp_1_0/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1098 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_651_413# 0.00fF
C1099 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_448_47# 0.00fF
C1100 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C1101 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_4/a_761_289# 0.00fF
C1102 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C1103 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_4/a_543_47# 0.00fF
C1104 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C1105 sky130_fd_sc_hd__nor3_2_3/B out 0.19fF
C1106 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C1107 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# SEL_CONV_TIME[2] 0.01fF
C1108 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__nor3_2_3/B 0.04fF
C1109 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C1110 sky130_fd_sc_hd__inv_1_48/A sky130_fd_sc_hd__nor3_2_3/B 0.41fF
C1111 sky130_fd_sc_hd__dfrtn_1_35/a_543_47# sky130_fd_sc_hd__dfrtn_1_36/a_1270_413# 0.00fF
C1112 sky130_fd_sc_hd__dfrtn_1_35/a_651_413# sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.00fF
C1113 sky130_fd_sc_hd__dfrtn_1_35/a_448_47# sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# 0.00fF
C1114 sky130_fd_sc_hd__dfrtn_1_37/a_639_47# sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# 0.00fF
C1115 sky130_fd_sc_hd__dfrtn_1_37/a_805_47# sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# 0.00fF
C1116 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# sky130_fd_sc_hd__dfrtn_1_39/a_1270_413# 0.00fF
C1117 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C1118 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C1119 sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C1120 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C1121 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_37/a_639_47# 0.00fF
C1122 sky130_fd_sc_hd__dfrtn_1_21/a_761_289# DOUT[2] 0.00fF
C1123 sky130_fd_sc_hd__dfrtn_1_9/a_805_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C1124 sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1125 sky130_fd_sc_hd__dfrtn_1_0/a_651_413# VDD 0.01fF
C1126 sky130_fd_sc_hd__dfrtn_1_35/a_543_47# VDD 0.06fF
C1127 sky130_fd_sc_hd__or2_2_0/B sky130_fd_sc_hd__or2_2_0/A 0.16fF
C1128 sky130_fd_sc_hd__nor3_2_2/A DOUT[15] 0.01fF
C1129 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__nor3_2_0/A 0.67fF
C1130 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__inv_1_15/A 0.01fF
C1131 sky130_fd_sc_hd__nor3_1_13/a_109_297# sky130_fd_sc_hd__dfrtn_1_8/a_543_47# 0.00fF
C1132 sky130_fd_sc_hd__dfrtn_1_3/a_651_413# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C1133 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# SEL_CONV_TIME[0] 0.01fF
C1134 sky130_fd_sc_hd__dfrtn_1_11/a_805_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C1135 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__inv_1_53/A 0.00fF
C1136 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# DOUT[19] 0.01fF
C1137 sky130_fd_sc_hd__nor3_1_2/a_193_297# DOUT[22] 0.00fF
C1138 sky130_fd_sc_hd__nor3_1_5/A DOUT[17] 0.00fF
C1139 sky130_fd_sc_hd__dfrtn_1_27/a_761_289# sky130_fd_sc_hd__or3_1_0/C 0.03fF
C1140 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# 0.00fF
C1141 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# SEL_CONV_TIME[0] 0.01fF
C1142 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C1143 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# VDD 0.14fF
C1144 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_14/a_448_47# -0.02fF
C1145 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C1146 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C1147 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_30/a_193_47# 0.00fF
C1148 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_24/a_543_47# 0.00fF
C1149 sky130_fd_sc_hd__dfrtn_1_20/a_1462_47# VDD 0.00fF
C1150 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C1151 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__inv_1_48/A 0.01fF
C1152 sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# RESET_COUNTERn 0.00fF
C1153 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_543_47# -0.00fF
C1154 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# -0.00fF
C1155 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# SLC_0/a_438_293# 0.00fF
C1156 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# RESET_COUNTERn 0.01fF
C1157 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C1158 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__inv_1_26/A 0.01fF
C1159 sky130_fd_sc_hd__dfrtn_1_9/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1160 CLK_REF sky130_fd_sc_hd__dfrtp_1_3/a_543_47# 0.01fF
C1161 DOUT[1] sky130_fd_sc_hd__dfrtn_1_36/a_1462_47# 0.00fF
C1162 DOUT[4] sky130_fd_sc_hd__dfrtn_1_8/a_1217_47# 0.00fF
C1163 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_2/a_448_47# 0.00fF
C1164 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_4/a_639_47# 0.00fF
C1165 sky130_fd_sc_hd__dfrtn_1_8/a_27_47# outb 0.00fF
C1166 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# -0.00fF
C1167 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_12/a_448_47# -0.00fF
C1168 sky130_fd_sc_hd__nand3b_1_0/a_53_93# SEL_CONV_TIME[1] 0.02fF
C1169 VDD sky130_fd_sc_hd__inv_1_44/A 0.46fF
C1170 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# -0.00fF
C1171 sky130_fd_sc_hd__dfrtn_1_16/a_639_47# DOUT[2] 0.00fF
C1172 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__dfrtn_1_13/a_193_47# 0.00fF
C1173 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_651_413# 0.00fF
C1174 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# 0.00fF
C1175 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# 0.00fF
C1176 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# sky130_fd_sc_hd__dfrtn_1_13/a_27_47# 0.00fF
C1177 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.01fF
C1178 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_12/a_27_47# 0.01fF
C1179 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# VIN 0.06fF
C1180 DOUT[9] sky130_fd_sc_hd__dfrtn_1_4/a_448_47# 0.00fF
C1181 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__inv_1_5/Y 0.18fF
C1182 sky130_fd_sc_hd__inv_1_31/Y RESET_COUNTERn 0.02fF
C1183 sky130_fd_sc_hd__nor3_1_17/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1184 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__dfrtp_1_0/a_448_47# -0.00fF
C1185 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__dfrtp_1_0/a_1108_47# -0.00fF
C1186 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1187 sky130_fd_sc_hd__o2111a_2_0/X DOUT[21] 0.00fF
C1188 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__inv_1_4/Y 0.01fF
C1189 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# SEL_CONV_TIME[0] 0.00fF
C1190 sky130_fd_sc_hd__dfrtn_1_37/a_639_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C1191 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_19/a_805_47# 0.00fF
C1192 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# VIN 0.01fF
C1193 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# 0.00fF
C1194 sky130_fd_sc_hd__mux4_2_0/X DOUT[21] 0.00fF
C1195 sky130_fd_sc_hd__dfrtn_1_34/a_543_47# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C1196 sky130_fd_sc_hd__nor3_1_2/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1197 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_20/a_1270_413# 0.00fF
C1198 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C1199 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_1217_47# -0.00fF
C1200 sky130_fd_sc_hd__nor3_1_11/a_193_297# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C1201 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# DOUT[21] 0.00fF
C1202 sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C1203 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# RESET_COUNTERn 0.01fF
C1204 sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C1205 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_11/a_805_47# 0.00fF
C1206 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# VDD 0.05fF
C1207 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# DOUT[7] 0.00fF
C1208 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# DOUT[20] 0.00fF
C1209 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# RESET_COUNTERn 0.01fF
C1210 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# sky130_fd_sc_hd__dfrtn_1_4/a_448_47# 0.00fF
C1211 sky130_fd_sc_hd__dfrtn_1_39/a_1217_47# SEL_CONV_TIME[2] 0.00fF
C1212 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_39/a_543_47# 0.01fF
C1213 sky130_fd_sc_hd__o311a_1_0/A3 sky130_fd_sc_hd__o2111a_2_0/X 0.08fF
C1214 SEL_CONV_TIME[1] sky130_fd_sc_hd__inv_1_43/A 0.11fF
C1215 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__inv_1_45/A 0.00fF
C1216 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_1270_413# 0.00fF
C1217 sky130_fd_sc_hd__dfrtn_1_33/a_1108_47# RESET_COUNTERn 0.00fF
C1218 DOUT[1] sky130_fd_sc_hd__dfrtn_1_32/a_1270_413# 0.00fF
C1219 sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# DOUT[19] 0.00fF
C1220 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__dfrtn_1_14/a_543_47# 0.00fF
C1221 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__dfrtn_1_14/a_761_289# 0.00fF
C1222 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_30/a_761_289# 0.00fF
C1223 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__mux4_2_0/a_872_316# 0.00fF
C1224 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__mux4_2_0/a_1060_369# 0.00fF
C1225 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__mux4_2_0/a_1279_413# 0.00fF
C1226 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C1227 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__o311a_1_0/A3 0.13fF
C1228 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1229 sky130_fd_sc_hd__dfrtn_1_30/a_805_47# RESET_COUNTERn 0.00fF
C1230 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_18/a_543_47# 0.00fF
C1231 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__inv_1_8/Y 0.01fF
C1232 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__inv_1_48/A 0.00fF
C1233 sky130_fd_sc_hd__nor3_1_11/a_193_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1234 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# 0.00fF
C1235 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C1236 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.00fF
C1237 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C1238 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__o311a_1_0/A3 0.01fF
C1239 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C1240 sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# SEL_CONV_TIME[0] 0.00fF
C1241 sky130_fd_sc_hd__mux4_2_0/a_397_47# SEL_CONV_TIME[1] -0.00fF
C1242 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# DOUT[19] 0.00fF
C1243 DOUT[19] DOUT[7] 0.02fF
C1244 sky130_fd_sc_hd__dfrtn_1_34/a_1462_47# SEL_CONV_TIME[0] 0.00fF
C1245 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C1246 sky130_fd_sc_hd__or3_1_0/a_111_297# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C1247 sky130_fd_sc_hd__dfrtn_1_17/a_761_289# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C1248 sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# VDD 0.00fF
C1249 sky130_fd_sc_hd__dfrtp_1_1/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1250 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C1251 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C1252 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# 0.00fF
C1253 sky130_fd_sc_hd__inv_1_39/A DOUT[14] 0.01fF
C1254 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C1255 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__inv_1_47/A 0.01fF
C1256 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C1257 sky130_fd_sc_hd__dfrtn_1_16/a_448_47# sky130_fd_sc_hd__inv_1_25/A 0.00fF
C1258 sky130_fd_sc_hd__dfrtp_1_0/a_805_47# SLC_0/a_264_22# 0.00fF
C1259 sky130_fd_sc_hd__dfrtp_1_0/a_1462_47# sky130_fd_sc_hd__inv_1_26/A 0.00fF
C1260 SLC_0/a_1235_416# out 0.00fF
C1261 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C1262 sky130_fd_sc_hd__dfrtn_1_38/a_543_47# RESET_COUNTERn 0.01fF
C1263 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# DOUT[18] 0.01fF
C1264 sky130_fd_sc_hd__nand3b_1_0/a_232_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C1265 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__nor3_1_5/a_193_297# 0.00fF
C1266 sky130_fd_sc_hd__dfrtn_1_14/a_543_47# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C1267 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C1268 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C1269 sky130_fd_sc_hd__dfrtn_1_17/a_1270_413# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C1270 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.00fF
C1271 sky130_fd_sc_hd__dfrtn_1_8/a_1217_47# outb 0.00fF
C1272 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1273 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_10/a_448_47# 0.00fF
C1274 sky130_fd_sc_hd__dfrtn_1_39/a_543_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C1275 sky130_fd_sc_hd__dfrtn_1_7/a_1462_47# VIN 0.00fF
C1276 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_12/a_1217_47# 0.00fF
C1277 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C1278 sky130_fd_sc_hd__mux4_2_0/a_872_316# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1279 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C1280 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C1281 sky130_fd_sc_hd__mux4_2_0/a_1279_413# VDD 0.00fF
C1282 sky130_fd_sc_hd__dfrtp_1_0/a_639_47# out 0.00fF
C1283 sky130_fd_sc_hd__nor3_1_10/a_193_297# sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# 0.00fF
C1284 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C1285 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# -0.00fF
C1286 out DOUT[0] 0.00fF
C1287 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C1288 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.00fF
C1289 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.03fF
C1290 sky130_fd_sc_hd__dfrtn_1_18/a_543_47# sky130_fd_sc_hd__inv_1_33/A 0.01fF
C1291 sky130_fd_sc_hd__dfrtn_1_27/a_651_413# SEL_CONV_TIME[1] 0.00fF
C1292 VDD sky130_fd_sc_hd__inv_1_32/A 1.67fF
C1293 sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# RESET_COUNTERn 0.02fF
C1294 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# 0.02fF
C1295 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C1296 sky130_fd_sc_hd__dfrtp_1_1/a_805_47# sky130_fd_sc_hd__nor3_2_1/a_27_297# 0.00fF
C1297 sky130_fd_sc_hd__dfrtn_1_33/a_448_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C1298 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C1299 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_543_47# 0.00fF
C1300 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.01fF
C1301 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__o211a_1_0/X 0.00fF
C1302 sky130_fd_sc_hd__dfrtn_1_35/a_639_47# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C1303 sky130_fd_sc_hd__dfrtn_1_16/a_1283_21# sky130_fd_sc_hd__nor3_2_3/A 0.02fF
C1304 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1305 sky130_fd_sc_hd__dfrtn_1_34/a_448_47# RESET_COUNTERn 0.00fF
C1306 sky130_fd_sc_hd__dfrtn_1_33/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1307 sky130_fd_sc_hd__dfrtn_1_11/a_1270_413# VDD 0.00fF
C1308 sky130_fd_sc_hd__dfrtn_1_35/a_1270_413# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C1309 sky130_fd_sc_hd__dfrtn_1_30/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1310 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_37/a_27_47# 0.00fF
C1311 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_37/a_193_47# 0.00fF
C1312 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_34/a_1270_413# 0.00fF
C1313 sky130_fd_sc_hd__dfrtn_1_8/a_448_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C1314 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_13/Y 0.08fF
C1315 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.01fF
C1316 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.01fF
C1317 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_35/a_543_47# 0.00fF
C1318 sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# DONE 0.00fF
C1319 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.00fF
C1320 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C1321 sky130_fd_sc_hd__inv_1_32/Y sky130_fd_sc_hd__inv_1_53/A 0.00fF
C1322 sky130_fd_sc_hd__dfrtn_1_28/a_1108_47# SEL_CONV_TIME[0] 0.00fF
C1323 sky130_fd_sc_hd__mux4_2_0/a_1064_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C1324 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__nand3b_1_0/a_316_47# 0.00fF
C1325 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C1326 DOUT[9] sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C1327 sky130_fd_sc_hd__dfrtn_1_38/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C1328 sky130_fd_sc_hd__dfrtn_1_27/a_448_47# VDD 0.01fF
C1329 sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1330 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C1331 sky130_fd_sc_hd__dfrtn_1_34/a_1217_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C1332 sky130_fd_sc_hd__inv_1_31/Y SEL_CONV_TIME[2] 0.00fF
C1333 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_18/a_448_47# 0.01fF
C1334 sky130_fd_sc_hd__nor3_1_18/a_193_297# VDD 0.00fF
C1335 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# RESET_COUNTERn 0.00fF
C1336 DOUT[4] sky130_fd_sc_hd__inv_1_38/A 0.15fF
C1337 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# 0.00fF
C1338 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C1339 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_448_47# -0.00fF
C1340 sky130_fd_sc_hd__dfrtn_1_36/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# -0.00fF
C1341 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C1342 sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C1343 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C1344 sky130_fd_sc_hd__o2111a_2_0/a_386_47# RESET_COUNTERn 0.00fF
C1345 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C1346 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C1347 sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C1348 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__a221oi_4_0/a_471_297# -0.00fF
C1349 sky130_fd_sc_hd__dfrtn_1_26/a_448_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C1350 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1351 sky130_fd_sc_hd__dfrtn_1_0/a_761_289# DOUT[18] 0.01fF
C1352 sky130_fd_sc_hd__dfrtn_1_26/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C1353 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# VDD 0.00fF
C1354 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C1355 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C1356 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# 0.00fF
C1357 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C1358 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__nor3_1_0/A 0.05fF
C1359 sky130_fd_sc_hd__nor3_1_19/a_193_297# RESET_COUNTERn 0.00fF
C1360 sky130_fd_sc_hd__dfrtp_1_3/a_1270_413# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C1361 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__o221ai_1_0/a_493_297# 0.00fF
C1362 sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C1363 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_27/a_761_289# 0.00fF
C1364 sky130_fd_sc_hd__dfrtn_1_12/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1365 sky130_fd_sc_hd__dfrtn_1_12/a_639_47# VDD 0.00fF
C1366 sky130_fd_sc_hd__a221oi_4_0/a_453_47# SEL_CONV_TIME[1] 0.00fF
C1367 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C1368 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_30/a_651_413# 0.00fF
C1369 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_1/a_543_47# 0.00fF
C1370 sky130_fd_sc_hd__dfrtn_1_28/a_1283_21# DOUT[21] 0.00fF
C1371 sky130_fd_sc_hd__dfrtn_1_33/a_1270_413# DOUT[23] 0.00fF
C1372 sky130_fd_sc_hd__dfrtn_1_14/a_761_289# sky130_fd_sc_hd__nor3_1_1/a_193_297# 0.00fF
C1373 sky130_fd_sc_hd__dfrtn_1_14/a_543_47# sky130_fd_sc_hd__nor3_1_1/a_109_297# 0.00fF
C1374 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C1375 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__inv_1_50/Y 0.08fF
C1376 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# DOUT[9] 0.00fF
C1377 sky130_fd_sc_hd__dfrtn_1_0/a_651_413# DOUT[5] 0.00fF
C1378 sky130_fd_sc_hd__dfrtn_1_11/a_805_47# DOUT[14] 0.00fF
C1379 sky130_fd_sc_hd__dfrtn_1_14/a_448_47# RESET_COUNTERn 0.00fF
C1380 sky130_fd_sc_hd__mux4_1_0/a_923_363# SEL_CONV_TIME[0] 0.00fF
C1381 sky130_fd_sc_hd__dfrtn_1_28/a_1270_413# sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C1382 DOUT[13] DONE 0.01fF
C1383 sky130_fd_sc_hd__dfrtn_1_42/a_1270_413# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C1384 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_34/a_639_47# 0.00fF
C1385 sky130_fd_sc_hd__or3b_2_0/a_27_47# SEL_CONV_TIME[1] 0.01fF
C1386 sky130_fd_sc_hd__inv_1_5/A RESET_COUNTERn 0.21fF
C1387 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C1388 sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# sky130_fd_sc_hd__dfrtp_1_3/a_651_413# 0.00fF
C1389 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__dfrtp_1_3/a_805_47# 0.00fF
C1390 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# sky130_fd_sc_hd__dfrtp_1_3/a_1217_47# 0.00fF
C1391 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C1392 sky130_fd_sc_hd__dfrtn_1_21/a_761_289# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C1393 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# VIN 0.00fF
C1394 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_51/Y 0.02fF
C1395 sky130_fd_sc_hd__or3_1_0/a_111_297# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C1396 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C1397 sky130_fd_sc_hd__dfrtn_1_36/a_639_47# sky130_fd_sc_hd__inv_1_40/A 0.00fF
C1398 sky130_fd_sc_hd__dfrtn_1_4/a_543_47# VIN 0.00fF
C1399 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# DOUT[22] 0.00fF
C1400 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C1401 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C1402 sky130_fd_sc_hd__dfrtn_1_40/a_1462_47# sky130_fd_sc_hd__dfrtn_1_37/a_27_47# 0.00fF
C1403 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__dfrtn_1_37/a_1270_413# 0.00fF
C1404 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_37/a_805_47# 0.00fF
C1405 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_37/a_639_47# 0.00fF
C1406 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__dfrtn_1_37/a_543_47# 0.00fF
C1407 sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# sky130_fd_sc_hd__dfrtn_1_37/a_193_47# 0.00fF
C1408 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__dfrtn_1_37/a_651_413# 0.00fF
C1409 sky130_fd_sc_hd__dfrtn_1_24/a_805_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C1410 DOUT[1] sky130_fd_sc_hd__dfrtn_1_23/a_27_47# 0.00fF
C1411 sky130_fd_sc_hd__a221oi_4_0/a_471_297# VDD 0.05fF
C1412 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C1413 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__dfrtn_1_2/a_651_413# 0.00fF
C1414 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# sky130_fd_sc_hd__dfrtn_1_2/a_761_289# 0.00fF
C1415 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C1416 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C1417 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# 0.00fF
C1418 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# 0.00fF
C1419 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# 0.00fF
C1420 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__dfrtn_1_2/a_805_47# 0.00fF
C1421 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_25/a_543_47# 0.00fF
C1422 sky130_fd_sc_hd__dfrtn_1_22/a_1283_21# sky130_fd_sc_hd__inv_1_39/A 0.01fF
C1423 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_24/a_651_413# -0.00fF
C1424 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C1425 sky130_fd_sc_hd__inv_1_13/Y DOUT[20] 0.00fF
C1426 sky130_fd_sc_hd__nor3_2_3/C SEL_CONV_TIME[1] 0.36fF
C1427 sky130_fd_sc_hd__dfrtn_1_42/a_448_47# DOUT[2] 0.00fF
C1428 sky130_fd_sc_hd__dfrtn_1_38/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1429 sky130_fd_sc_hd__or3b_2_0/a_176_21# VDD 0.09fF
C1430 DOUT[1] sky130_fd_sc_hd__dfrtn_1_22/a_805_47# 0.00fF
C1431 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# SEL_CONV_TIME[1] 0.02fF
C1432 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_543_47# -0.00fF
C1433 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_34/a_543_47# 0.01fF
C1434 DOUT[13] sky130_fd_sc_hd__nor3_2_3/B 0.07fF
C1435 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# RESET_COUNTERn 0.01fF
C1436 DOUT[4] sky130_fd_sc_hd__o221ai_1_0/a_493_297# 0.00fF
C1437 sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C1438 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_41/a_448_47# 0.01fF
C1439 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_19/a_543_47# 0.01fF
C1440 sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# DOUT[23] 0.00fF
C1441 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# DOUT[14] 0.00fF
C1442 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# DOUT[19] 0.01fF
C1443 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__inv_1_8/A 0.06fF
C1444 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__dfrtn_1_15/a_543_47# 0.00fF
C1445 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# 0.00fF
C1446 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_639_47# 0.00fF
C1447 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C1448 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__dfrtn_1_15/a_761_289# 0.00fF
C1449 sky130_fd_sc_hd__dfrtn_1_25/a_651_413# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C1450 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1451 sky130_fd_sc_hd__dfrtn_1_5/a_805_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C1452 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# 0.00fF
C1453 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C1454 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_805_47# 0.00fF
C1455 sky130_fd_sc_hd__dfrtn_1_5/a_805_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C1456 sky130_fd_sc_hd__dfrtn_1_17/a_761_289# VDD 0.04fF
C1457 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C1458 sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C1459 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__inv_1_54/Y 0.00fF
C1460 sky130_fd_sc_hd__dfrtn_1_14/a_651_413# sky130_fd_sc_hd__nor3_1_0/a_193_297# 0.00fF
C1461 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C1462 sky130_fd_sc_hd__dfrtn_1_36/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1463 sky130_fd_sc_hd__dfrtn_1_36/a_639_47# VDD 0.00fF
C1464 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_805_47# 0.00fF
C1465 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# 0.00fF
C1466 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__nor3_1_19/Y 0.01fF
C1467 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__o2111a_2_0/a_80_21# 0.00fF
C1468 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__o2111a_2_0/a_80_21# 0.00fF
C1469 sky130_fd_sc_hd__nor3_2_3/a_281_297# sky130_fd_sc_hd__dfrtn_1_42/a_543_47# 0.00fF
C1470 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# 0.00fF
C1471 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C1472 DOUT[11] DOUT[22] 0.01fF
C1473 sky130_fd_sc_hd__inv_1_17/A DOUT[12] 0.00fF
C1474 sky130_fd_sc_hd__dfrtn_1_0/a_1217_47# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C1475 sky130_fd_sc_hd__dfrtn_1_3/a_761_289# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C1476 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C1477 sky130_fd_sc_hd__o2111a_2_0/a_386_47# SEL_CONV_TIME[3] 0.00fF
C1478 sky130_fd_sc_hd__o311a_1_0/a_266_297# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C1479 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C1480 sky130_fd_sc_hd__dfrtn_1_28/a_805_47# RESET_COUNTERn 0.00fF
C1481 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# VDD 0.23fF
C1482 sky130_fd_sc_hd__dfrtn_1_39/a_1217_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C1483 sky130_fd_sc_hd__mux4_2_0/a_288_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C1484 sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C1485 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__nor3_1_1/a_109_297# 0.00fF
C1486 sky130_fd_sc_hd__mux4_2_0/a_27_47# SEL_CONV_TIME[0] 0.01fF
C1487 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_11/a_1270_413# 0.00fF
C1488 sky130_fd_sc_hd__dfrtn_1_0/a_543_47# RESET_COUNTERn 0.00fF
C1489 sky130_fd_sc_hd__inv_1_54/A DOUT[2] 0.01fF
C1490 sky130_fd_sc_hd__dfrtn_1_3/a_651_413# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C1491 sky130_fd_sc_hd__inv_1_43/Y sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C1492 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__o221ai_1_0/a_493_297# 0.00fF
C1493 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C1494 sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C1495 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C1496 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C1497 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# 0.00fF
C1498 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# 0.00fF
C1499 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_39/a_27_47# 0.00fF
C1500 sky130_fd_sc_hd__inv_1_49/Y DOUT[4] 0.01fF
C1501 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_30/a_543_47# 0.00fF
C1502 sky130_fd_sc_hd__nor3_1_3/a_193_297# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C1503 sky130_fd_sc_hd__nor3_1_4/a_109_297# VDD 0.00fF
C1504 sky130_fd_sc_hd__nor3_1_5/a_193_297# RESET_COUNTERn 0.00fF
C1505 outb sky130_fd_sc_hd__inv_1_11/Y 0.09fF
C1506 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C1507 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C1508 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__dfrtn_1_9/a_448_47# 0.00fF
C1509 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C1510 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_19/a_761_289# 0.00fF
C1511 sky130_fd_sc_hd__dfrtn_1_0/a_761_289# DOUT[22] 0.00fF
C1512 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__inv_1_31/A 0.11fF
C1513 sky130_fd_sc_hd__dfrtn_1_21/a_651_413# sky130_fd_sc_hd__inv_1_35/Y 0.00fF
C1514 sky130_fd_sc_hd__dfrtn_1_32/a_639_47# sky130_fd_sc_hd__inv_1_9/A 0.00fF
C1515 sky130_fd_sc_hd__dfrtn_1_20/a_1270_413# RESET_COUNTERn 0.00fF
C1516 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# SEL_CONV_TIME[0] 0.00fF
C1517 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_38/a_761_289# 0.00fF
C1518 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__o221ai_1_0/a_295_297# 0.00fF
C1519 sky130_fd_sc_hd__dfrtp_1_2/a_448_47# sky130_fd_sc_hd__inv_1_29/Y 0.00fF
C1520 DOUT[1] sky130_fd_sc_hd__dfrtn_1_23/a_1217_47# 0.00fF
C1521 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C1522 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# 0.00fF
C1523 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C1524 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_18/a_543_47# 0.00fF
C1525 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_448_47# 0.00fF
C1526 sky130_fd_sc_hd__dfrtn_1_18/a_639_47# DOUT[2] 0.00fF
C1527 sky130_fd_sc_hd__o2111a_2_0/a_386_47# SEL_CONV_TIME[2] 0.00fF
C1528 CLK_REF sky130_fd_sc_hd__dfrtp_1_1/D 0.02fF
C1529 sky130_fd_sc_hd__dfrtn_1_42/a_543_47# sky130_fd_sc_hd__inv_1_25/A 0.01fF
C1530 sky130_fd_sc_hd__dfrtn_1_32/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C1531 sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# VDD 0.07fF
C1532 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C1533 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# sky130_fd_sc_hd__inv_1_6/Y 0.11fF
C1534 sky130_fd_sc_hd__nor3_2_1/a_27_297# VDD 0.05fF
C1535 sky130_fd_sc_hd__nand3b_1_0/a_232_47# SEL_CONV_TIME[0] 0.00fF
C1536 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# DOUT[11] 0.00fF
C1537 sky130_fd_sc_hd__dfrtn_1_4/a_543_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C1538 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_38/a_448_47# 0.00fF
C1539 sky130_fd_sc_hd__dfrtn_1_36/a_543_47# sky130_fd_sc_hd__inv_1_52/Y 0.01fF
C1540 en DOUT[19] 0.06fF
C1541 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C1542 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__or2_2_0/A 0.24fF
C1543 DOUT[1] RESET_COUNTERn 0.06fF
C1544 sky130_fd_sc_hd__mux4_1_0/a_27_47# RESET_COUNTERn 0.01fF
C1545 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# 0.00fF
C1546 sky130_fd_sc_hd__nor3_2_1/A RESET_COUNTERn 0.03fF
C1547 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C1548 sky130_fd_sc_hd__o211a_1_0/a_215_47# RESET_COUNTERn 0.00fF
C1549 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.00fF
C1550 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_639_47# 0.00fF
C1551 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_31/a_805_47# 0.00fF
C1552 sky130_fd_sc_hd__or3b_2_0/a_472_297# sky130_fd_sc_hd__dfrtn_1_31/a_651_413# 0.00fF
C1553 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C1554 sky130_fd_sc_hd__o211a_1_0/a_79_21# lc_out 0.02fF
C1555 sky130_fd_sc_hd__dfrtn_1_42/a_193_47# sky130_fd_sc_hd__nor3_2_3/A 0.02fF
C1556 sky130_fd_sc_hd__dfrtn_1_28/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1557 sky130_fd_sc_hd__dfrtn_1_21/a_1462_47# DOUT[2] 0.00fF
C1558 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C1559 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C1560 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# DOUT[9] 0.00fF
C1561 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# VDD 0.04fF
C1562 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__inv_1_33/A 0.01fF
C1563 sky130_fd_sc_hd__dfrtn_1_22/a_639_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C1564 sky130_fd_sc_hd__inv_1_27/Y sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1565 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__conb_1_0/LO 0.00fF
C1566 DOUT[4] sky130_fd_sc_hd__inv_1_0/Y 0.01fF
C1567 DOUT[4] sky130_fd_sc_hd__dfrtn_1_30/a_543_47# 0.00fF
C1568 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__dfrtn_1_30/a_448_47# -0.00fF
C1569 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# -0.00fF
C1570 sky130_fd_sc_hd__nand3b_1_0/a_53_93# DOUT[21] 0.00fF
C1571 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_639_47# 0.00fF
C1572 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_448_47# 0.00fF
C1573 sky130_fd_sc_hd__nor3_1_9/a_109_297# DOUT[11] 0.00fF
C1574 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C1575 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C1576 sky130_fd_sc_hd__or2_2_0/B RESET_COUNTERn 0.45fF
C1577 sky130_fd_sc_hd__nor3_1_11/a_109_297# sky130_fd_sc_hd__dfrtn_1_7/a_448_47# 0.00fF
C1578 sky130_fd_sc_hd__dfrtn_1_19/a_27_47# sky130_fd_sc_hd__inv_1_28/A 0.48fF
C1579 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfrtn_1_41/a_448_47# -0.02fF
C1580 sky130_fd_sc_hd__dfrtn_1_31/a_1217_47# VDD 0.00fF
C1581 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C1582 sky130_fd_sc_hd__mux4_2_0/a_1064_47# SEL_CONV_TIME[0] 0.00fF
C1583 sky130_fd_sc_hd__dfrtn_1_38/a_448_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C1584 sky130_fd_sc_hd__dfrtn_1_28/a_448_47# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C1585 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C1586 VDD sky130_fd_sc_hd__inv_1_9/Y 0.30fF
C1587 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C1588 sky130_fd_sc_hd__dfrtn_1_35/a_805_47# RESET_COUNTERn 0.00fF
C1589 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# sky130_fd_sc_hd__dfrtn_1_31/a_639_47# -0.00fF
C1590 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_805_47# -0.00fF
C1591 sky130_fd_sc_hd__nor3_1_11/a_109_297# DOUT[8] 0.00fF
C1592 sky130_fd_sc_hd__nor3_1_11/a_193_297# DOUT[7] 0.00fF
C1593 CLK_REF sky130_fd_sc_hd__dfrtn_1_21/a_651_413# 0.00fF
C1594 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# DOUT[3] 0.00fF
C1595 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_14/a_543_47# 0.00fF
C1596 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# RESET_COUNTERn 0.00fF
C1597 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__dfrtn_1_25/a_27_47# 0.00fF
C1598 sky130_fd_sc_hd__dfrtn_1_4/a_639_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C1599 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C1600 sky130_fd_sc_hd__dfrtp_1_3/a_543_47# sky130_fd_sc_hd__dfrtn_1_17/a_543_47# 0.00fF
C1601 sky130_fd_sc_hd__dfrtp_1_3/a_761_289# sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# 0.00fF
C1602 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# 0.00fF
C1603 sky130_fd_sc_hd__dfrtp_1_3/a_448_47# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C1604 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_448_47# 0.00fF
C1605 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# DOUT[18] 0.00fF
C1606 sky130_fd_sc_hd__dfrtn_1_40/a_1462_47# sky130_fd_sc_hd__inv_1_31/A 0.00fF
C1607 sky130_fd_sc_hd__inv_1_31/Y sky130_fd_sc_hd__inv_1_53/A 0.00fF
C1608 sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C1609 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtp_1_2/a_193_47# -0.00fF
C1610 sky130_fd_sc_hd__dfrtn_1_12/a_761_289# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C1611 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C1612 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__dfrtn_1_18/a_1462_47# 0.00fF
C1613 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_18/a_1217_47# 0.00fF
C1614 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C1615 sky130_fd_sc_hd__dfrtn_1_4/a_761_289# sky130_fd_sc_hd__inv_1_7/A 0.01fF
C1616 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__dfrtn_1_29/a_448_47# 0.00fF
C1617 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__dfrtn_1_29/a_543_47# 0.00fF
C1618 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# 0.00fF
C1619 sky130_fd_sc_hd__dfrtn_1_10/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1620 sky130_fd_sc_hd__o211a_1_0/a_79_21# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C1621 sky130_fd_sc_hd__dfrtp_1_3/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1622 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C1623 sky130_fd_sc_hd__dfrtp_1_3/a_1108_47# VDD 0.07fF
C1624 sky130_fd_sc_hd__inv_1_43/A DOUT[21] 0.00fF
C1625 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# SEL_CONV_TIME[1] 0.00fF
C1626 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_21/a_193_47# 0.01fF
C1627 sky130_fd_sc_hd__dfrtp_1_3/a_1462_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C1628 sky130_fd_sc_hd__inv_1_36/A sky130_fd_sc_hd__inv_1_39/Y 0.01fF
C1629 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C1630 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# 0.00fF
C1631 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# 0.00fF
C1632 sky130_fd_sc_hd__dfrtn_1_27/a_1270_413# SEL_CONV_TIME[0] 0.00fF
C1633 sky130_fd_sc_hd__mux4_2_0/a_600_345# RESET_COUNTERn 0.00fF
C1634 sky130_fd_sc_hd__dfrtn_1_23/a_805_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C1635 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/D 0.00fF
C1636 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_36/a_639_47# 0.00fF
C1637 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__inv_1_47/A 0.00fF
C1638 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_543_47# -0.00fF
C1639 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_761_289# -0.00fF
C1640 sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C1641 sky130_fd_sc_hd__dfrtn_1_4/a_805_47# DOUT[11] 0.00fF
C1642 sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# RESET_COUNTERn 0.02fF
C1643 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__dfrtn_1_33/a_651_413# -0.00fF
C1644 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# sky130_fd_sc_hd__dfrtn_1_33/a_448_47# -0.00fF
C1645 sky130_fd_sc_hd__dfrtn_1_0/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1646 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1647 sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# DOUT[9] 0.00fF
C1648 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# DOUT[19] 0.00fF
C1649 sky130_fd_sc_hd__dfrtn_1_35/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1650 sky130_fd_sc_hd__nor3_2_0/a_27_297# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C1651 sky130_fd_sc_hd__nor3_1_15/a_109_297# VDD 0.00fF
C1652 sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C1653 sky130_fd_sc_hd__dfrtn_1_40/a_1462_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C1654 sky130_fd_sc_hd__dfrtn_1_41/a_639_47# RESET_COUNTERn 0.00fF
C1655 sky130_fd_sc_hd__dfrtn_1_0/a_1462_47# sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# 0.00fF
C1656 sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# sky130_fd_sc_hd__dfrtn_1_3/a_1462_47# 0.00fF
C1657 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_34/a_805_47# 0.00fF
C1658 sky130_fd_sc_hd__nor3_2_1/a_27_297# sky130_fd_sc_hd__o211a_1_0/X 0.00fF
C1659 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C1660 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# VDD 0.01fF
C1661 DOUT[4] outb 0.02fF
C1662 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C1663 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1664 sky130_fd_sc_hd__dfrtn_1_3/a_805_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C1665 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__o211a_1_1/a_510_47# 0.00fF
C1666 sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.01fF
C1667 sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C1668 HEADER_1/a_508_138# VDD 0.04fF
C1669 sky130_fd_sc_hd__dfrtn_1_32/a_805_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C1670 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# sky130_fd_sc_hd__o211a_1_1/X 0.00fF
C1671 sky130_fd_sc_hd__dfrtn_1_23/a_761_289# sky130_fd_sc_hd__dfrtn_1_36/a_543_47# 0.00fF
C1672 sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.01fF
C1673 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C1674 sky130_fd_sc_hd__dfrtn_1_27/a_651_413# DOUT[21] 0.00fF
C1675 sky130_fd_sc_hd__dfrtn_1_27/a_761_289# RESET_COUNTERn 0.01fF
C1676 sky130_fd_sc_hd__dfrtn_1_38/a_543_47# sky130_fd_sc_hd__inv_1_53/A 0.01fF
C1677 sky130_fd_sc_hd__dfrtn_1_35/a_543_47# sky130_fd_sc_hd__inv_1_38/A 0.01fF
C1678 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C1679 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# 0.00fF
C1680 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__dfrtn_1_25/a_448_47# 0.00fF
C1681 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_25/a_651_413# 0.00fF
C1682 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__dfrtn_1_25/a_193_47# 0.00fF
C1683 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_25/a_805_47# 0.00fF
C1684 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# 0.00fF
C1685 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__inv_1_49/A 0.02fF
C1686 sky130_fd_sc_hd__nor3_2_0/a_27_297# sky130_fd_sc_hd__dfrtn_1_12/a_27_47# 0.00fF
C1687 sky130_fd_sc_hd__o311a_1_0/a_368_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1688 sky130_fd_sc_hd__dfrtn_1_38/a_193_47# DOUT[2] 0.00fF
C1689 sky130_fd_sc_hd__inv_1_21/Y VIN 0.10fF
C1690 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C1691 sky130_fd_sc_hd__dfrtn_1_37/a_1270_413# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C1692 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# sky130_fd_sc_hd__mux4_2_0/a_372_413# 0.00fF
C1693 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# sky130_fd_sc_hd__mux4_2_0/a_600_345# 0.00fF
C1694 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__mux4_2_0/a_872_316# 0.00fF
C1695 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# sky130_fd_sc_hd__mux4_2_0/a_193_47# 0.00fF
C1696 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# sky130_fd_sc_hd__mux4_2_0/a_193_369# 0.00fF
C1697 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C1698 sky130_fd_sc_hd__dfrtn_1_10/a_1283_21# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C1699 sky130_fd_sc_hd__mux4_2_0/a_372_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1700 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C1701 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# sky130_fd_sc_hd__nor3_1_2/a_109_297# 0.00fF
C1702 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# sky130_fd_sc_hd__nor3_1_2/a_193_297# 0.00fF
C1703 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C1704 sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C1705 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# SEL_CONV_TIME[0] 0.01fF
C1706 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# RESET_COUNTERn 0.02fF
C1707 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# sky130_fd_sc_hd__inv_1_13/Y 0.01fF
C1708 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C1709 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__nor3_1_4/A 1.10fF
C1710 sky130_fd_sc_hd__nor3_1_10/a_193_297# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C1711 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C1712 sky130_fd_sc_hd__dfrtn_1_33/a_543_47# sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# 0.00fF
C1713 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_651_413# 0.00fF
C1714 DOUT[12] DOUT[21] 0.00fF
C1715 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C1716 sky130_fd_sc_hd__dfrtn_1_34/a_1270_413# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C1717 sky130_fd_sc_hd__dfrtn_1_22/a_651_413# VDD 0.01fF
C1718 sky130_fd_sc_hd__dfrtn_1_22/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1719 sky130_fd_sc_hd__dfrtn_1_11/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1720 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# RESET_COUNTERn 0.00fF
C1721 sky130_fd_sc_hd__dfrtn_1_39/a_193_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C1722 sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# 0.00fF
C1723 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_543_47# -0.00fF
C1724 sky130_fd_sc_hd__dfrtn_1_38/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_761_289# -0.00fF
C1725 DOUT[1] sky130_fd_sc_hd__dfrtn_1_42/a_1108_47# 0.00fF
C1726 sky130_fd_sc_hd__dfrtn_1_41/a_805_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C1727 sky130_fd_sc_hd__dfrtn_1_28/a_639_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C1728 sky130_fd_sc_hd__nor3_1_20/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1729 sky130_fd_sc_hd__nor3_1_4/a_109_297# DOUT[3] 0.00fF
C1730 sky130_fd_sc_hd__dfrtn_1_41/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1731 DOUT[4] sky130_fd_sc_hd__dfrtn_1_34/a_805_47# 0.00fF
C1732 sky130_fd_sc_hd__dfrtn_1_26/a_543_47# DOUT[2] 0.00fF
C1733 sky130_fd_sc_hd__or3b_2_0/a_388_297# SEL_CONV_TIME[0] 0.00fF
C1734 sky130_fd_sc_hd__dfrtn_1_18/a_193_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C1735 sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# sky130_fd_sc_hd__dfrtp_1_1/D 0.00fF
C1736 DOUT[19] VIN 3.73fF
C1737 sky130_fd_sc_hd__dfrtn_1_23/a_1270_413# sky130_fd_sc_hd__inv_1_40/A 0.00fF
C1738 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__dfrtp_1_1/a_543_47# 0.00fF
C1739 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# sky130_fd_sc_hd__dfrtp_1_1/a_27_47# 0.00fF
C1740 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/a_761_289# 0.00fF
C1741 sky130_fd_sc_hd__nor3_1_4/a_109_297# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C1742 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.00fF
C1743 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C1744 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.00fF
C1745 sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C1746 sky130_fd_sc_hd__o311a_1_0/a_585_47# SEL_CONV_TIME[3] 0.00fF
C1747 sky130_fd_sc_hd__dfrtn_1_8/a_1108_47# sky130_fd_sc_hd__inv_1_9/A 0.01fF
C1748 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_10/a_805_47# 0.00fF
C1749 sky130_fd_sc_hd__dfrtp_1_1/a_805_47# DOUT[23] 0.00fF
C1750 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# DOUT[19] 0.00fF
C1751 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C1752 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C1753 sky130_fd_sc_hd__dfrtn_1_27/a_543_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C1754 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C1755 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C1756 sky130_fd_sc_hd__dfrtn_1_8/a_805_47# DOUT[12] 0.00fF
C1757 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_2/Y 0.01fF
C1758 sky130_fd_sc_hd__dfrtn_1_3/a_651_413# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C1759 sky130_fd_sc_hd__nor3_2_1/A SLC_0/a_264_22# 0.01fF
C1760 sky130_fd_sc_hd__inv_1_15/A sky130_fd_sc_hd__nor3_2_3/B 0.40fF
C1761 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C1762 sky130_fd_sc_hd__mux4_2_0/a_600_345# SEL_CONV_TIME[3] 0.01fF
C1763 sky130_fd_sc_hd__dfrtn_1_16/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C1764 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.03fF
C1765 sky130_fd_sc_hd__dfrtn_1_16/a_1108_47# VDD 0.07fF
C1766 SLC_0/a_264_22# sky130_fd_sc_hd__o211a_1_0/a_215_47# 0.00fF
C1767 sky130_fd_sc_hd__dfrtn_1_8/a_193_47# VDD 0.09fF
C1768 sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C1769 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C1770 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C1771 sky130_fd_sc_hd__a221oi_4_0/a_453_47# DOUT[21] 0.00fF
C1772 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__inv_1_47/A 0.01fF
C1773 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__inv_1_9/Y 0.01fF
C1774 CLK_REF sky130_fd_sc_hd__dfrtn_1_19/a_805_47# 0.00fF
C1775 sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C1776 sky130_fd_sc_hd__dfrtn_1_21/a_805_47# sky130_fd_sc_hd__inv_1_35/A 0.00fF
C1777 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1778 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_20/a_543_47# 0.01fF
C1779 sky130_fd_sc_hd__dfrtn_1_18/a_639_47# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C1780 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__dfrtn_1_29/a_639_47# 0.00fF
C1781 sky130_fd_sc_hd__dfrtn_1_31/a_761_289# SEL_CONV_TIME[0] 0.01fF
C1782 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# DOUT[2] 0.00fF
C1783 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# -0.00fF
C1784 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C1785 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C1786 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_34/a_805_47# 0.00fF
C1787 sky130_fd_sc_hd__dfrtp_1_0/a_639_47# sky130_fd_sc_hd__o211a_1_0/a_79_21# 0.00fF
C1788 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C1789 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_651_413# -0.00fF
C1790 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__dfrtn_1_26/a_448_47# -0.00fF
C1791 sky130_fd_sc_hd__o211a_1_0/a_79_21# DOUT[0] 0.00fF
C1792 sky130_fd_sc_hd__o211a_1_0/a_297_297# out 0.00fF
C1793 sky130_fd_sc_hd__nor3_1_12/a_109_297# DOUT[21] 0.00fF
C1794 DOUT[9] sky130_fd_sc_hd__inv_1_13/A 0.00fF
C1795 sky130_fd_sc_hd__o311a_1_0/a_585_47# SEL_CONV_TIME[2] 0.00fF
C1796 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1797 SLC_0/a_264_22# sky130_fd_sc_hd__or2_2_0/B 0.01fF
C1798 sky130_fd_sc_hd__dfrtn_1_9/a_761_289# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C1799 sky130_fd_sc_hd__mux4_2_0/a_600_345# SEL_CONV_TIME[2] 0.00fF
C1800 sky130_fd_sc_hd__dfrtn_1_23/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1801 sky130_fd_sc_hd__inv_1_39/A sky130_fd_sc_hd__inv_1_40/Y 0.07fF
C1802 sky130_fd_sc_hd__dfrtn_1_9/a_639_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C1803 sky130_fd_sc_hd__inv_1_50/A SEL_CONV_TIME[1] 0.15fF
C1804 sky130_fd_sc_hd__dfrtn_1_23/a_1270_413# VDD 0.00fF
C1805 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1806 sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C1807 DOUT[13] sky130_fd_sc_hd__dfrtn_1_30/a_639_47# 0.00fF
C1808 sky130_fd_sc_hd__dfrtn_1_38/a_1462_47# DOUT[2] 0.00fF
C1809 sky130_fd_sc_hd__dfrtn_1_37/a_1462_47# sky130_fd_sc_hd__mux4_2_0/a_872_316# 0.00fF
C1810 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_639_47# 0.00fF
C1811 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C1812 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_38/a_543_47# 0.00fF
C1813 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C1814 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__o311a_1_0/A3 0.01fF
C1815 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_3/a_193_47# 0.00fF
C1816 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1817 sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# VDD 0.08fF
C1818 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# DOUT[14] 0.14fF
C1819 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__inv_1_29/Y 0.00fF
C1820 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__inv_1_13/A 0.01fF
C1821 sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# RESET_COUNTERn 0.03fF
C1822 sky130_fd_sc_hd__dfrtn_1_36/a_805_47# DOUT[21] 0.00fF
C1823 sky130_fd_sc_hd__dfrtn_1_37/a_805_47# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C1824 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C1825 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C1826 sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C1827 sky130_fd_sc_hd__o311a_1_0/a_368_297# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C1828 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# VDD 0.00fF
C1829 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1830 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C1831 sky130_fd_sc_hd__inv_1_44/Y sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C1832 sky130_fd_sc_hd__nor3_2_3/C DOUT[21] 0.33fF
C1833 VDD DOUT[6] 1.20fF
C1834 sky130_fd_sc_hd__dfrtn_1_20/a_651_413# sky130_fd_sc_hd__dfrtn_1_21/a_1462_47# 0.00fF
C1835 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__o311a_1_0/A3 0.07fF
C1836 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__dfrtn_1_25/a_805_47# 0.00fF
C1837 sky130_fd_sc_hd__inv_1_42/A sky130_fd_sc_hd__or3_1_0/C 0.01fF
C1838 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C1839 sky130_fd_sc_hd__dfrtn_1_18/a_1462_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C1840 sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# RESET_COUNTERn 0.03fF
C1841 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C1842 sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# DOUT[23] 0.00fF
C1843 sky130_fd_sc_hd__dfrtp_1_0/a_805_47# sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# 0.00fF
C1844 sky130_fd_sc_hd__dfrtp_1_0/a_639_47# sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# 0.00fF
C1845 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# 0.00fF
C1846 sky130_fd_sc_hd__dfrtp_1_0/a_761_289# sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# 0.00fF
C1847 sky130_fd_sc_hd__or3_1_0/a_183_297# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C1848 sky130_fd_sc_hd__nor3_1_18/a_109_297# DOUT[23] 0.00fF
C1849 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# 0.00fF
C1850 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# SEL_CONV_TIME[1] 0.00fF
C1851 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# 0.00fF
C1852 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# sky130_fd_sc_hd__dfrtn_1_27/a_543_47# 0.00fF
C1853 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# 0.00fF
C1854 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_448_47# 0.00fF
C1855 sky130_fd_sc_hd__dfrtn_1_25/a_448_47# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C1856 sky130_fd_sc_hd__or2b_1_0/X sky130_fd_sc_hd__inv_1_42/A 0.00fF
C1857 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C1858 sky130_fd_sc_hd__nor3_1_4/a_109_297# DOUT[20] 0.00fF
C1859 sky130_fd_sc_hd__o2111a_2_0/a_458_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C1860 sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# sky130_fd_sc_hd__inv_1_37/A 0.03fF
C1861 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C1862 sky130_fd_sc_hd__dfrtn_1_27/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1863 sky130_fd_sc_hd__dfrtn_1_8/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1864 sky130_fd_sc_hd__dfrtn_1_8/a_1462_47# VDD 0.00fF
C1865 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__o311a_1_0/A3 0.10fF
C1866 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C1867 sky130_fd_sc_hd__dfrtn_1_34/a_651_413# sky130_fd_sc_hd__inv_1_49/A 0.01fF
C1868 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# -0.00fF
C1869 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C1870 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C1871 DOUT[13] sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# 0.00fF
C1872 sky130_fd_sc_hd__dfrtn_1_23/a_761_289# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C1873 sky130_fd_sc_hd__dfrtn_1_32/a_193_47# RESET_COUNTERn 0.00fF
C1874 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__dfrtn_1_34/a_543_47# 0.00fF
C1875 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C1876 sky130_fd_sc_hd__dfrtn_1_8/a_27_47# sky130_fd_sc_hd__inv_1_9/Y 0.24fF
C1877 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# CLK_REF 0.02fF
C1878 sky130_fd_sc_hd__o311a_1_0/a_266_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C1879 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__dfrtn_1_22/a_761_289# -0.00fF
C1880 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__inv_1_1/Y 0.00fF
C1881 sky130_fd_sc_hd__dfrtn_1_36/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1882 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_15/a_193_47# 0.00fF
C1883 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C1884 sky130_fd_sc_hd__inv_1_6/A sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C1885 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C1886 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C1887 sky130_fd_sc_hd__dfrtn_1_5/a_805_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C1888 sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# sky130_fd_sc_hd__inv_1_44/A 0.02fF
C1889 sky130_fd_sc_hd__dfrtn_1_7/a_448_47# DOUT[14] 0.00fF
C1890 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# VDD -0.20fF
C1891 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C1892 sky130_fd_sc_hd__dfrtn_1_25/a_1270_413# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C1893 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.13fF
C1894 sky130_fd_sc_hd__nor3_2_0/a_281_297# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C1895 outb sky130_fd_sc_hd__nor3_2_3/A 0.03fF
C1896 sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# sky130_fd_sc_hd__inv_1_32/A 0.01fF
C1897 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__mux4_2_0/a_1060_369# 0.00fF
C1898 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_3/a_1462_47# 0.00fF
C1899 sky130_fd_sc_hd__dfrtn_1_17/a_639_47# RESET_COUNTERn 0.00fF
C1900 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# DOUT[14] 0.00fF
C1901 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__o2111a_2_0/a_674_297# -0.00fF
C1902 sky130_fd_sc_hd__dfrtn_1_41/a_1270_413# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C1903 DOUT[8] DOUT[14] 0.50fF
C1904 sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C1905 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1906 sky130_fd_sc_hd__inv_1_29/A VDD 0.27fF
C1907 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C1908 sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# sky130_fd_sc_hd__inv_1_32/A 0.01fF
C1909 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_1270_413# 0.00fF
C1910 sky130_fd_sc_hd__or3b_2_0/B VDD 0.91fF
C1911 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C1912 sky130_fd_sc_hd__dfrtn_1_0/a_651_413# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C1913 sky130_fd_sc_hd__dfrtn_1_19/a_193_47# sky130_fd_sc_hd__inv_1_34/Y 0.08fF
C1914 DOUT[4] sky130_fd_sc_hd__dfrtn_1_35/a_543_47# 0.00fF
C1915 sky130_fd_sc_hd__dfrtn_1_11/a_1270_413# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C1916 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C1917 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_805_47# 0.00fF
C1918 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_639_47# 0.00fF
C1919 sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__inv_1_41/Y 0.17fF
C1920 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C1921 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__inv_1_35/A 0.05fF
C1922 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C1923 sky130_fd_sc_hd__dfrtn_1_31/a_651_413# RESET_COUNTERn 0.00fF
C1924 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C1925 sky130_fd_sc_hd__nand3b_1_0/Y RESET_COUNTERn 0.00fF
C1926 sky130_fd_sc_hd__dfrtn_1_20/a_1270_413# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C1927 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_4/a_1270_413# 0.00fF
C1928 sky130_fd_sc_hd__inv_1_27/Y DOUT[2] 0.02fF
C1929 DOUT[1] sky130_fd_sc_hd__nor3_2_2/A 0.01fF
C1930 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_12/a_761_289# 0.00fF
C1931 sky130_fd_sc_hd__dfrtn_1_9/a_651_413# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C1932 sky130_fd_sc_hd__or2_2_0/a_39_297# sky130_fd_sc_hd__dfrtn_1_19/a_651_413# 0.00fF
C1933 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# SEL_CONV_TIME[1] 0.00fF
C1934 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C1935 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# 0.00fF
C1936 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_8/a_193_47# 0.01fF
C1937 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_31/a_639_47# 0.00fF
C1938 sky130_fd_sc_hd__dfrtn_1_33/a_1462_47# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C1939 sky130_fd_sc_hd__dfrtn_1_20/a_448_47# DOUT[2] 0.00fF
C1940 sky130_fd_sc_hd__dfrtn_1_22/a_543_47# sky130_fd_sc_hd__dfrtn_1_23/a_27_47# 0.00fF
C1941 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__dfrtn_1_23/a_543_47# 0.00fF
C1942 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_21/a_543_47# 0.01fF
C1943 sky130_fd_sc_hd__dfrtn_1_31/a_1108_47# DONE 0.00fF
C1944 sky130_fd_sc_hd__mux4_2_0/a_1060_369# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C1945 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_21/a_27_47# 0.05fF
C1946 sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C1947 sky130_fd_sc_hd__dfrtn_1_38/a_761_289# sky130_fd_sc_hd__inv_1_27/Y 0.00fF
C1948 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# 0.00fF
C1949 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C1950 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__dfrtp_1_1/D 0.20fF
C1951 outb sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C1952 sky130_fd_sc_hd__dfrtn_1_29/a_805_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C1953 sky130_fd_sc_hd__dfrtn_1_32/a_1462_47# RESET_COUNTERn 0.00fF
C1954 sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# SEL_CONV_TIME[0] 0.00fF
C1955 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_33/a_1108_47# 0.00fF
C1956 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__dfrtn_1_33/a_27_47# 0.00fF
C1957 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# 0.00fF
C1958 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_33/a_1270_413# 0.00fF
C1959 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__dfrtn_1_33/a_448_47# 0.00fF
C1960 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# RESET_COUNTERn 0.01fF
C1961 sky130_fd_sc_hd__dfrtn_1_8/a_1217_47# sky130_fd_sc_hd__inv_1_9/Y 0.00fF
C1962 sky130_fd_sc_hd__dfrtn_1_28/a_805_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C1963 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.00fF
C1964 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C1965 sky130_fd_sc_hd__dfrtn_1_17/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C1966 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# outb 0.00fF
C1967 VDD DOUT[23] 4.82fF
C1968 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_23/a_1270_413# 0.00fF
C1969 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# VDD 0.08fF
C1970 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C1971 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C1972 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_27_47# 0.00fF
C1973 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C1974 sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# VDD 0.00fF
C1975 sky130_fd_sc_hd__dfrtn_1_12/a_651_413# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C1976 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_17/a_1462_47# 0.00fF
C1977 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__inv_1_46/Y 0.00fF
C1978 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__inv_1_35/Y 0.02fF
C1979 sky130_fd_sc_hd__dfrtn_1_3/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C1980 sky130_fd_sc_hd__dfrtn_1_3/a_805_47# VDD 0.00fF
C1981 sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C1982 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# 0.00fF
C1983 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__dfrtp_1_2/a_193_47# 0.00fF
C1984 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_2/a_448_47# 0.00fF
C1985 sky130_fd_sc_hd__dfrtp_1_1/a_448_47# sky130_fd_sc_hd__dfrtp_1_2/a_27_47# 0.00fF
C1986 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__dfrtp_1_2/a_543_47# 0.00fF
C1987 sky130_fd_sc_hd__dfrtn_1_34/a_448_47# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C1988 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C1989 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C1990 sky130_fd_sc_hd__nor3_2_1/a_281_297# sky130_fd_sc_hd__dfrtp_1_1/D 0.01fF
C1991 sky130_fd_sc_hd__nor3_1_2/a_193_297# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C1992 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C1993 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C1994 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C1995 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# 0.00fF
C1996 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_639_47# 0.00fF
C1997 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C1998 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C1999 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# RESET_COUNTERn 0.00fF
C2000 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__inv_1_44/A 0.02fF
C2001 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C2002 sky130_fd_sc_hd__dfrtn_1_42/a_761_289# VDD 0.03fF
C2003 sky130_fd_sc_hd__dfrtn_1_19/a_1462_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C2004 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# DOUT[21] 0.00fF
C2005 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# RESET_COUNTERn 0.03fF
C2006 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__inv_1_8/A 0.02fF
C2007 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_36/a_761_289# 0.00fF
C2008 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# -0.00fF
C2009 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# sky130_fd_sc_hd__dfrtn_1_23/a_543_47# -0.00fF
C2010 DOUT[11] sky130_fd_sc_hd__inv_1_8/A 0.00fF
C2011 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C2012 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# VDD 0.04fF
C2013 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C2014 sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.03fF
C2015 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# DOUT[11] 0.00fF
C2016 sky130_fd_sc_hd__dfrtn_1_4/a_448_47# VDD 0.01fF
C2017 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# 0.00fF
C2018 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# 0.00fF
C2019 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C2020 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_761_289# 0.00fF
C2021 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__dfrtn_1_26/a_805_47# 0.00fF
C2022 sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.00fF
C2023 sky130_fd_sc_hd__nor3_1_0/A DOUT[18] 0.04fF
C2024 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__inv_1_31/A 0.00fF
C2025 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__nor3_1_1/a_193_297# 0.00fF
C2026 sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# DOUT[3] 0.02fF
C2027 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# 0.00fF
C2028 sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C2029 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_8/a_1462_47# 0.00fF
C2030 sky130_fd_sc_hd__dfrtn_1_19/a_639_47# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C2031 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# sky130_fd_sc_hd__dfrtn_1_16/a_639_47# -0.00fF
C2032 sky130_fd_sc_hd__dfrtn_1_8/a_27_47# sky130_fd_sc_hd__dfrtn_1_8/a_193_47# -0.08fF
C2033 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# DOUT[3] 0.00fF
C2034 DOUT[6] DOUT[3] 0.00fF
C2035 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C2036 DOUT[9] sky130_fd_sc_hd__inv_1_3/A 0.00fF
C2037 sky130_fd_sc_hd__nand3b_1_0/Y SEL_CONV_TIME[3] 0.16fF
C2038 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C2039 sky130_fd_sc_hd__o311a_1_0/a_585_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C2040 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__dfrtn_1_7/a_193_47# 0.01fF
C2041 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_761_289# 0.00fF
C2042 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# sky130_fd_sc_hd__dfrtn_1_7/a_27_47# 0.00fF
C2043 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C2044 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__nor3_1_4/a_193_297# 0.00fF
C2045 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# 0.02fF
C2046 sky130_fd_sc_hd__or2b_1_0/a_301_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2047 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__dfrtn_1_16/a_1270_413# 0.00fF
C2048 sky130_fd_sc_hd__nor3_2_2/a_281_297# sky130_fd_sc_hd__dfrtn_1_16/a_651_413# 0.00fF
C2049 sky130_fd_sc_hd__mux4_2_0/a_600_345# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C2050 sky130_fd_sc_hd__dfrtn_1_28/a_193_47# sky130_fd_sc_hd__dfrtn_1_28/a_1108_47# -0.00fF
C2051 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__dfrtn_1_28/a_448_47# -0.00fF
C2052 sky130_fd_sc_hd__dfrtp_1_0/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2053 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__nor3_2_3/B 0.04fF
C2054 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C2055 sky130_fd_sc_hd__dfrtp_1_0/a_1283_21# VDD 0.11fF
C2056 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C2057 sky130_fd_sc_hd__inv_1_2/A DOUT[6] 0.01fF
C2058 sky130_fd_sc_hd__dfrtp_1_1/a_805_47# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C2059 sky130_fd_sc_hd__dfrtp_1_3/a_1462_47# RESET_COUNTERn 0.00fF
C2060 sky130_fd_sc_hd__dfrtp_1_1/a_639_47# sky130_fd_sc_hd__o211a_1_1/a_215_47# 0.00fF
C2061 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C2062 sky130_fd_sc_hd__dfrtn_1_22/a_543_47# RESET_COUNTERn 0.00fF
C2063 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C2064 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_448_47# 0.00fF
C2065 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C2066 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C2067 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C2068 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C2069 sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# VDD 0.08fF
C2070 CLK_REF sky130_fd_sc_hd__dfrtn_1_20/a_27_47# 0.01fF
C2071 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2072 sky130_fd_sc_hd__dfrtn_1_25/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2073 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C2074 sky130_fd_sc_hd__dfrtn_1_25/a_1462_47# VDD 0.00fF
C2075 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C2076 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_10/a_193_47# -0.16fF
C2077 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# sky130_fd_sc_hd__dfrtn_1_3/a_27_47# 0.00fF
C2078 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__dfrtn_1_3/a_193_47# 0.00fF
C2079 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_3/a_805_47# 0.00fF
C2080 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__dfrtn_1_3/a_639_47# 0.00fF
C2081 sky130_fd_sc_hd__nor3_1_11/a_193_297# VIN 0.00fF
C2082 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C2083 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C2084 sky130_fd_sc_hd__o221ai_1_0/a_213_123# SEL_CONV_TIME[1] 0.00fF
C2085 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__inv_1_33/A 0.05fF
C2086 sky130_fd_sc_hd__inv_1_31/A VDD 0.53fF
C2087 sky130_fd_sc_hd__nor3_2_3/a_281_297# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C2088 sky130_fd_sc_hd__nand3b_1_0/Y SEL_CONV_TIME[2] 0.01fF
C2089 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C2090 sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# VDD 0.09fF
C2091 DOUT[9] sky130_fd_sc_hd__nor3_2_3/C 0.40fF
C2092 sky130_fd_sc_hd__dfrtn_1_20/a_1217_47# sky130_fd_sc_hd__inv_1_35/Y 0.00fF
C2093 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__o221ai_1_0/a_295_297# 0.00fF
C2094 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__o221ai_1_0/a_493_297# 0.00fF
C2095 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# sky130_fd_sc_hd__inv_1_5/Y 0.03fF
C2096 sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C2097 sky130_fd_sc_hd__dfrtn_1_41/a_651_413# DOUT[2] 0.00fF
C2098 sky130_fd_sc_hd__dfrtp_1_1/a_805_47# sky130_fd_sc_hd__dfrtp_1_2/a_651_413# 0.00fF
C2099 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__dfrtp_1_2/a_805_47# 0.00fF
C2100 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C2101 sky130_fd_sc_hd__dfrtn_1_17/a_193_47# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C2102 sky130_fd_sc_hd__dfrtn_1_17/a_761_289# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C2103 sky130_fd_sc_hd__dfrtn_1_24/a_805_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C2104 sky130_fd_sc_hd__dfrtn_1_42/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2105 sky130_fd_sc_hd__dfrtn_1_16/a_193_47# RESET_COUNTERn -0.02fF
C2106 sky130_fd_sc_hd__dfrtn_1_8/a_761_289# DOUT[21] 0.00fF
C2107 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# DOUT[14] 0.00fF
C2108 sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C2109 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C2110 VDD sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.05fF
C2111 sky130_fd_sc_hd__nor3_1_6/a_193_297# RESET_COUNTERn 0.00fF
C2112 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_20/a_761_289# -0.00fF
C2113 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_651_413# 0.00fF
C2114 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C2115 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C2116 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C2117 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__mux4_2_0/a_1279_413# 0.00fF
C2118 sky130_fd_sc_hd__dfrtn_1_10/a_1462_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C2119 sky130_fd_sc_hd__dfrtn_1_41/a_639_47# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C2120 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C2121 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.01fF
C2122 sky130_fd_sc_hd__dfrtn_1_41/a_1270_413# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C2123 sky130_fd_sc_hd__dfrtn_1_41/a_651_413# sky130_fd_sc_hd__dfrtn_1_38/a_761_289# 0.00fF
C2124 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# sky130_fd_sc_hd__dfrtn_1_38/a_448_47# 0.00fF
C2125 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# sky130_fd_sc_hd__dfrtn_1_38/a_651_413# 0.00fF
C2126 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_639_47# 0.00fF
C2127 sky130_fd_sc_hd__dfrtn_1_19/a_193_47# VDD 0.08fF
C2128 DOUT[9] sky130_fd_sc_hd__nor3_1_4/a_193_297# 0.00fF
C2129 sky130_fd_sc_hd__dfrtp_1_3/a_1283_21# DOUT[23] 0.00fF
C2130 sky130_fd_sc_hd__nor3_2_2/a_27_297# RESET_COUNTERn 0.01fF
C2131 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2132 sky130_fd_sc_hd__inv_1_28/Y sky130_fd_sc_hd__o211a_1_1/X 0.00fF
C2133 DOUT[23] sky130_fd_sc_hd__o211a_1_0/X 0.00fF
C2134 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__or2b_1_0/a_27_53# 0.00fF
C2135 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C2136 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# 0.00fF
C2137 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_1/a_448_47# 0.00fF
C2138 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_1/a_193_47# 0.00fF
C2139 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_1/a_27_47# 0.00fF
C2140 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_1/a_651_413# 0.00fF
C2141 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C2142 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# 0.00fF
C2143 sky130_fd_sc_hd__o221ai_1_0/a_295_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2144 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__mux4_2_0/a_1060_369# 0.00fF
C2145 sky130_fd_sc_hd__o221ai_1_0/a_109_47# VDD 0.01fF
C2146 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.07fF
C2147 sky130_fd_sc_hd__dfrtn_1_24/a_448_47# SEL_CONV_TIME[1] 0.00fF
C2148 sky130_fd_sc_hd__inv_1_37/A sky130_fd_sc_hd__inv_1_36/A 0.01fF
C2149 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# sky130_fd_sc_hd__o221ai_1_0/a_295_297# 0.00fF
C2150 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__o221ai_1_0/a_493_297# 0.00fF
C2151 sky130_fd_sc_hd__dfrtp_1_3/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2152 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# sky130_fd_sc_hd__dfrtn_1_7/a_448_47# -0.00fF
C2153 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_651_413# -0.00fF
C2154 VDD sky130_fd_sc_hd__inv_1_33/A 3.77fF
C2155 sky130_fd_sc_hd__dfrtn_1_16/a_639_47# DOUT[15] 0.00fF
C2156 sky130_fd_sc_hd__dfrtn_1_33/a_1270_413# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C2157 sky130_fd_sc_hd__nor3_1_4/a_109_297# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C2158 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C2159 sky130_fd_sc_hd__nor3_1_1/a_109_297# DOUT[18] 0.00fF
C2160 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# RESET_COUNTERn 0.03fF
C2161 sky130_fd_sc_hd__dfrtn_1_23/a_639_47# DOUT[21] 0.00fF
C2162 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2163 sky130_fd_sc_hd__dfrtn_1_26/a_448_47# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C2164 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__or3b_2_0/a_176_21# 0.00fF
C2165 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__dfrtn_1_26/a_448_47# 0.00fF
C2166 sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C2167 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__dfrtn_1_26/a_651_413# 0.00fF
C2168 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__dfrtn_1_7/a_1462_47# 0.00fF
C2169 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# sky130_fd_sc_hd__dfrtn_1_7/a_193_47# 0.00fF
C2170 DOUT[4] sky130_fd_sc_hd__dfrtn_1_12/a_639_47# 0.00fF
C2171 sky130_fd_sc_hd__dfrtn_1_10/a_1283_21# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C2172 sky130_fd_sc_hd__dfrtn_1_12/a_639_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C2173 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# DOUT[7] 0.00fF
C2174 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# RESET_COUNTERn 0.02fF
C2175 sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# DOUT[20] 0.00fF
C2176 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# DOUT[8] 0.00fF
C2177 sky130_fd_sc_hd__dfrtn_1_7/a_543_47# DOUT[6] 0.00fF
C2178 sky130_fd_sc_hd__dfrtn_1_21/a_543_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C2179 sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C2180 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_0/a_543_47# -0.00fF
C2181 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# sky130_fd_sc_hd__dfrtn_1_0/a_761_289# -0.00fF
C2182 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# DOUT[6] 0.00fF
C2183 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# RESET_COUNTERn 0.00fF
C2184 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# DOUT[20] 0.00fF
C2185 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# DOUT[7] 0.00fF
C2186 DOUT[20] DOUT[6] 9.73fF
C2187 DOUT[22] sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C2188 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C2189 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__mux4_1_0/a_277_47# -0.00fF
C2190 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_32/a_639_47# 0.00fF
C2191 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C2192 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C2193 sky130_fd_sc_hd__dfrtn_1_27/a_761_289# sky130_fd_sc_hd__inv_1_42/Y 0.01fF
C2194 sky130_fd_sc_hd__dfrtn_1_26/a_543_47# sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.00fF
C2195 sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C2196 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2197 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__o311a_1_0/a_266_47# 0.00fF
C2198 sky130_fd_sc_hd__o2111a_2_0/a_458_47# sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.00fF
C2199 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# VDD 0.07fF
C2200 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C2201 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C2202 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# VDD 0.15fF
C2203 sky130_fd_sc_hd__dfrtn_1_11/a_1270_413# outb 0.00fF
C2204 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__or3_1_0/C 0.30fF
C2205 sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2206 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# SEL_CONV_TIME[0] 0.00fF
C2207 sky130_fd_sc_hd__inv_1_43/Y SEL_CONV_TIME[0] 0.27fF
C2208 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__dfrtn_1_3/a_543_47# 0.00fF
C2209 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_31/a_27_47# 0.07fF
C2210 sky130_fd_sc_hd__nor3_1_3/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2211 sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# DOUT[14] 0.00fF
C2212 sky130_fd_sc_hd__or3b_2_0/X SEL_CONV_TIME[1] 0.01fF
C2213 sky130_fd_sc_hd__inv_1_34/Y sky130_fd_sc_hd__inv_1_35/Y 0.00fF
C2214 sky130_fd_sc_hd__inv_1_9/Y sky130_fd_sc_hd__inv_1_11/Y 0.01fF
C2215 outb sky130_fd_sc_hd__inv_1_19/A 0.01fF
C2216 sky130_fd_sc_hd__dfrtn_1_17/a_1462_47# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C2217 sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# sky130_fd_sc_hd__dfrtn_1_19/a_639_47# 0.00fF
C2218 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# SEL_CONV_TIME[1] 0.00fF
C2219 sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C2220 sky130_fd_sc_hd__dfrtn_1_16/a_1462_47# RESET_COUNTERn 0.00fF
C2221 sky130_fd_sc_hd__dfrtn_1_8/a_1270_413# RESET_COUNTERn 0.00fF
C2222 sky130_fd_sc_hd__dfrtp_1_0/a_1283_21# sky130_fd_sc_hd__o211a_1_0/X 0.00fF
C2223 sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2224 sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# SEL_CONV_TIME[1] 0.03fF
C2225 sky130_fd_sc_hd__dfrtn_1_20/a_448_47# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C2226 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_21/a_639_47# 0.00fF
C2227 sky130_fd_sc_hd__dfrtn_1_32/a_651_413# sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C2228 DOUT[4] sky130_fd_sc_hd__or3b_2_0/a_176_21# 0.00fF
C2229 sky130_fd_sc_hd__dfrtn_1_23/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2230 sky130_fd_sc_hd__dfrtn_1_19/a_1462_47# VDD 0.00fF
C2231 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2232 sky130_fd_sc_hd__or3b_2_0/a_472_297# sky130_fd_sc_hd__dfrtn_1_30/a_27_47# 0.00fF
C2233 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__o311a_1_0/A3 0.15fF
C2234 sky130_fd_sc_hd__dfrtn_1_24/a_651_413# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C2235 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C2236 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# VDD -0.23fF
C2237 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__or2_2_0/A 0.01fF
C2238 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C2239 sky130_fd_sc_hd__nor3_1_10/a_193_297# sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# 0.00fF
C2240 sky130_fd_sc_hd__dfrtn_1_34/a_651_413# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C2241 sky130_fd_sc_hd__dfrtn_1_22/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2242 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C2243 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# 0.00fF
C2244 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__inv_1_47/Y 0.01fF
C2245 sky130_fd_sc_hd__o311a_1_0/a_81_21# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C2246 sky130_fd_sc_hd__inv_1_48/Y sky130_fd_sc_hd__nor3_2_3/B 0.03fF
C2247 sky130_fd_sc_hd__dfrtn_1_7/a_1217_47# RESET_COUNTERn 0.00fF
C2248 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_29/a_805_47# 0.00fF
C2249 sky130_fd_sc_hd__dfrtn_1_30/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2250 sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# VDD 0.09fF
C2251 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# DOUT[3] 0.00fF
C2252 sky130_fd_sc_hd__dfrtn_1_4/a_448_47# DOUT[3] 0.00fF
C2253 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__a221oi_4_0/a_27_297# 0.00fF
C2254 sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C2255 sky130_fd_sc_hd__dfrtn_1_16/a_1283_21# DOUT[23] 0.00fF
C2256 DOUT[4] sky130_fd_sc_hd__dfrtn_1_31/a_27_47# 0.00fF
C2257 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__inv_1_48/A 0.01fF
C2258 sky130_fd_sc_hd__dfrtn_1_30/a_543_47# sky130_fd_sc_hd__dfrtn_1_31/a_27_47# 0.00fF
C2259 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_543_47# 0.00fF
C2260 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# DOUT[14] 0.00fF
C2261 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__or3_1_0/X 0.01fF
C2262 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__dfrtn_1_35/a_448_47# -0.00fF
C2263 sky130_fd_sc_hd__nor3_1_1/a_193_297# RESET_COUNTERn 0.00fF
C2264 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# sky130_fd_sc_hd__inv_1_15/A 0.01fF
C2265 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__inv_1_2/A 0.01fF
C2266 sky130_fd_sc_hd__dfrtp_1_1/a_805_47# CLK_REF 0.00fF
C2267 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C2268 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C2269 sky130_fd_sc_hd__dfrtn_1_4/a_448_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C2270 sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# DOUT[17] 0.00fF
C2271 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__mux4_1_0/a_1478_413# -0.00fF
C2272 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_834_97# -0.00fF
C2273 sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# sky130_fd_sc_hd__dfrtn_1_27/a_543_47# 0.00fF
C2274 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# SEL_CONV_TIME[1] 0.01fF
C2275 sky130_fd_sc_hd__o211a_1_1/a_215_47# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C2276 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__dfrtn_1_17/a_761_289# 0.00fF
C2277 sky130_fd_sc_hd__o211a_1_1/a_297_297# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C2278 sky130_fd_sc_hd__dfrtn_1_16/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2279 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# SEL_CONV_TIME[0] 0.00fF
C2280 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2281 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# VDD -0.00fF
C2282 sky130_fd_sc_hd__dfrtn_1_8/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2283 sky130_fd_sc_hd__o211a_1_0/a_79_21# sky130_fd_sc_hd__o211a_1_0/a_297_297# -0.00fF
C2284 sky130_fd_sc_hd__dfrtn_1_36/a_448_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C2285 CLK_REF sky130_fd_sc_hd__inv_1_34/Y 0.01fF
C2286 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C2287 sky130_fd_sc_hd__or2_2_0/X VDD 0.16fF
C2288 sky130_fd_sc_hd__nor3_1_1/a_109_297# DOUT[22] 0.00fF
C2289 sky130_fd_sc_hd__nand3b_1_0/a_316_47# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C2290 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C2291 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__nor3_1_3/a_109_297# 0.00fF
C2292 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_543_47# 0.00fF
C2293 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# sky130_fd_sc_hd__dfrtn_1_11/a_193_47# 0.00fF
C2294 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_11/a_761_289# 0.00fF
C2295 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__dfrtn_1_11/a_27_47# 0.00fF
C2296 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C2297 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C2298 sky130_fd_sc_hd__o211a_1_1/a_297_297# VDD 0.00fF
C2299 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# 0.00fF
C2300 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_12/a_651_413# 0.00fF
C2301 DOUT[4] sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# 0.00fF
C2302 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__inv_1_54/A 0.20fF
C2303 VDD sky130_fd_sc_hd__o2111a_2_0/X 0.18fF
C2304 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__dfrtn_1_40/a_193_47# 0.00fF
C2305 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__dfrtn_1_40/a_543_47# 0.00fF
C2306 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C2307 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_17/a_543_47# 0.00fF
C2308 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# 0.01fF
C2309 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C2310 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_651_413# 0.00fF
C2311 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_14/a_651_413# 0.00fF
C2312 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__dfrtn_1_14/a_761_289# 0.00fF
C2313 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# 0.00fF
C2314 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# 0.00fF
C2315 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C2316 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_14/a_761_289# 0.00fF
C2317 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__or3_1_0/C 0.01fF
C2318 sky130_fd_sc_hd__inv_1_13/A sky130_fd_sc_hd__inv_1_8/Y 0.02fF
C2319 sky130_fd_sc_hd__mux4_2_0/X VDD 0.25fF
C2320 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C2321 sky130_fd_sc_hd__dfrtn_1_20/a_639_47# sky130_fd_sc_hd__dfrtn_1_21/a_27_47# 0.00fF
C2322 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C2323 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# DOUT[14] 0.01fF
C2324 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# VDD -0.18fF
C2325 sky130_fd_sc_hd__dfrtn_1_10/a_1283_21# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C2326 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# VDD 0.01fF
C2327 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__dfrtn_1_30/a_27_47# 0.00fF
C2328 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# sky130_fd_sc_hd__o221ai_1_0/a_295_297# 0.00fF
C2329 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C2330 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C2331 sky130_fd_sc_hd__dfrtn_1_7/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2332 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C2333 DOUT[11] sky130_fd_sc_hd__inv_1_15/A 0.02fF
C2334 SLC_0/a_919_243# sky130_fd_sc_hd__dfrtn_1_16/a_27_47# 0.00fF
C2335 sky130_fd_sc_hd__dfrtn_1_16/a_543_47# sky130_fd_sc_hd__inv_1_26/A 0.00fF
C2336 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2337 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# VDD 0.00fF
C2338 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# DOUT[21] 0.00fF
C2339 sky130_fd_sc_hd__dfrtn_1_12/a_651_413# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C2340 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_6/a_543_47# 0.00fF
C2341 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# RESET_COUNTERn 0.01fF
C2342 sky130_fd_sc_hd__dfrtn_1_32/a_761_289# sky130_fd_sc_hd__inv_1_36/A 0.02fF
C2343 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C2344 sky130_fd_sc_hd__dfrtn_1_9/a_761_289# DOUT[3] 0.00fF
C2345 DOUT[9] sky130_fd_sc_hd__dfrtn_1_6/a_27_47# 0.00fF
C2346 sky130_fd_sc_hd__dfrtn_1_33/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2347 sky130_fd_sc_hd__dfrtn_1_33/a_805_47# VDD 0.00fF
C2348 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# RESET_COUNTERn 0.01fF
C2349 sky130_fd_sc_hd__dfrtn_1_31/a_639_47# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C2350 sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__or3_1_0/C 0.01fF
C2351 lc_out sky130_fd_sc_hd__nor3_2_3/B 0.26fF
C2352 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C2353 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C2354 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__inv_1_53/A 0.00fF
C2355 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# HEADER_0/a_508_138# 0.00fF
C2356 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2357 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# VDD 0.06fF
C2358 sky130_fd_sc_hd__dfrtn_1_20/a_805_47# sky130_fd_sc_hd__inv_1_35/A 0.00fF
C2359 sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C2360 sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C2361 sky130_fd_sc_hd__dfrtn_1_21/a_543_47# VDD 0.05fF
C2362 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C2363 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C2364 sky130_fd_sc_hd__inv_1_37/A sky130_fd_sc_hd__inv_1_7/A 0.00fF
C2365 sky130_fd_sc_hd__nor3_1_19/Y sky130_fd_sc_hd__inv_1_41/Y 0.12fF
C2366 sky130_fd_sc_hd__nand3b_1_1/Y sky130_fd_sc_hd__inv_1_48/A 0.00fF
C2367 DONE sky130_fd_sc_hd__nor3_2_3/B 0.09fF
C2368 sky130_fd_sc_hd__inv_1_50/Y SEL_CONV_TIME[0] 0.06fF
C2369 sky130_fd_sc_hd__or2b_1_0/X sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C2370 sky130_fd_sc_hd__dfrtn_1_0/a_761_289# sky130_fd_sc_hd__inv_1_15/A 0.01fF
C2371 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C2372 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# HEADER_0/a_508_138# 0.00fF
C2373 sky130_fd_sc_hd__inv_1_42/A RESET_COUNTERn 0.21fF
C2374 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# sky130_fd_sc_hd__or2_2_0/B 0.03fF
C2375 DOUT[13] sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.00fF
C2376 sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# DOUT[17] 0.00fF
C2377 sky130_fd_sc_hd__dfrtn_1_34/a_1462_47# SEL_CONV_TIME[1] 0.00fF
C2378 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# DOUT[20] 0.00fF
C2379 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# DOUT[8] 0.00fF
C2380 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# DOUT[7] 0.00fF
C2381 sky130_fd_sc_hd__dfrtn_1_24/a_805_47# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C2382 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C2383 sky130_fd_sc_hd__dfrtn_1_24/a_651_413# sky130_fd_sc_hd__dfrtn_1_29/a_543_47# 0.00fF
C2384 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_29/a_639_47# 0.00fF
C2385 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# sky130_fd_sc_hd__dfrtn_1_29/a_651_413# 0.00fF
C2386 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_805_47# 0.00fF
C2387 sky130_fd_sc_hd__dfrtn_1_17/a_761_289# sky130_fd_sc_hd__inv_1_28/A 0.01fF
C2388 sky130_fd_sc_hd__dfrtn_1_8/a_193_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C2389 DOUT[13] sky130_fd_sc_hd__inv_1_9/A 0.00fF
C2390 sky130_fd_sc_hd__nand3b_1_1/a_316_47# RESET_COUNTERn 0.00fF
C2391 sky130_fd_sc_hd__dfrtn_1_4/a_761_289# RESET_COUNTERn 0.01fF
C2392 sky130_fd_sc_hd__or3_1_0/a_183_297# RESET_COUNTERn 0.00fF
C2393 sky130_fd_sc_hd__dfrtn_1_38/a_1270_413# VDD 0.00fF
C2394 sky130_fd_sc_hd__dfrtn_1_33/a_448_47# sky130_fd_sc_hd__inv_1_45/A 0.01fF
C2395 sky130_fd_sc_hd__nor3_1_5/a_109_297# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C2396 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__dfrtn_1_11/a_1217_47# 0.00fF
C2397 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__dfrtn_1_11/a_1270_413# 0.00fF
C2398 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# sky130_fd_sc_hd__dfrtn_1_11/a_1462_47# 0.00fF
C2399 sky130_fd_sc_hd__dfrtn_1_10/a_639_47# sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# 0.00fF
C2400 sky130_fd_sc_hd__dfrtn_1_10/a_805_47# sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# 0.00fF
C2401 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# sky130_fd_sc_hd__dfrtn_1_11/a_651_413# 0.00fF
C2402 sky130_fd_sc_hd__inv_1_9/A sky130_fd_sc_hd__inv_1_8/A 0.00fF
C2403 sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C2404 sky130_fd_sc_hd__dfrtn_1_42/a_448_47# DOUT[15] 0.00fF
C2405 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/a_805_47# -0.00fF
C2406 sky130_fd_sc_hd__dfrtn_1_7/a_805_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C2407 HEADER_2/a_508_138# VIN 0.03fF
C2408 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__dfrtn_1_40/a_1462_47# 0.00fF
C2409 sky130_fd_sc_hd__dfrtn_1_12/a_651_413# sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# 0.00fF
C2410 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# VDD 0.15fF
C2411 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# 0.00fF
C2412 VDD sky130_fd_sc_hd__inv_1_35/Y 0.32fF
C2413 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C2414 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_37/a_805_47# -0.00fF
C2415 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# 0.00fF
C2416 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# 0.01fF
C2417 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__dfrtn_1_0/a_193_47# 0.01fF
C2418 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# sky130_fd_sc_hd__dfrtn_1_0/a_27_47# 0.00fF
C2419 sky130_fd_sc_hd__or2_2_0/a_39_297# sky130_fd_sc_hd__or2_2_0/B 0.01fF
C2420 sky130_fd_sc_hd__dfrtn_1_28/a_1217_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C2421 sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2422 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2423 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__inv_1_45/A 0.01fF
C2424 sky130_fd_sc_hd__dfrtn_1_26/a_805_47# VDD 0.00fF
C2425 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# DOUT[3] 0.00fF
C2426 sky130_fd_sc_hd__inv_1_17/A VIN 0.10fF
C2427 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# RESET_COUNTERn 0.01fF
C2428 sky130_fd_sc_hd__inv_1_48/A sky130_fd_sc_hd__inv_1_51/Y 0.05fF
C2429 sky130_fd_sc_hd__nor3_1_10/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2430 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__dfrtn_1_41/a_543_47# -0.00fF
C2431 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C2432 sky130_fd_sc_hd__dfrtn_1_34/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2433 sky130_fd_sc_hd__dfrtn_1_34/a_1217_47# VDD 0.00fF
C2434 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C2435 sky130_fd_sc_hd__nor3_1_11/a_109_297# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C2436 sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2437 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# 0.00fF
C2438 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# 0.00fF
C2439 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_8/a_1108_47# 0.01fF
C2440 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.01fF
C2441 sky130_fd_sc_hd__dfrtn_1_23/a_805_47# sky130_fd_sc_hd__inv_1_40/Y 0.00fF
C2442 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C2443 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__inv_1_42/Y 0.03fF
C2444 SLC_0/a_919_243# DOUT[15] 0.00fF
C2445 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_3/a_651_413# -0.00fF
C2446 sky130_fd_sc_hd__dfrtn_1_41/a_805_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C2447 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__inv_1_2/A 0.02fF
C2448 sky130_fd_sc_hd__dfrtn_1_21/a_639_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C2449 sky130_fd_sc_hd__dfrtn_1_39/a_193_47# RESET_COUNTERn 0.00fF
C2450 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__inv_1_7/A 0.00fF
C2451 sky130_fd_sc_hd__nor3_1_19/Y sky130_fd_sc_hd__inv_1_49/A 0.00fF
C2452 DOUT[13] sky130_fd_sc_hd__dfrtn_1_32/a_27_47# 0.00fF
C2453 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_21/a_1217_47# 0.00fF
C2454 sky130_fd_sc_hd__dfrtn_1_25/a_1270_413# RESET_COUNTERn 0.00fF
C2455 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__inv_1_54/A 0.01fF
C2456 sky130_fd_sc_hd__dfrtp_1_3/a_1283_21# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C2457 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C2458 sky130_fd_sc_hd__nor3_1_15/a_109_297# DOUT[4] 0.00fF
C2459 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C2460 sky130_fd_sc_hd__dfrtn_1_18/a_193_47# RESET_COUNTERn 0.00fF
C2461 DOUT[9] DOUT[7] 0.01fF
C2462 sky130_fd_sc_hd__dfrtp_1_0/a_1270_413# DOUT[15] 0.00fF
C2463 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_26/a_448_47# 0.01fF
C2464 DOUT[15] out 0.41fF
C2465 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C2466 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2467 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C2468 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__inv_1_43/A 0.01fF
C2469 sky130_fd_sc_hd__dfrtn_1_7/a_1217_47# HEADER_0/a_508_138# 0.00fF
C2470 sky130_fd_sc_hd__dfrtn_1_28/a_1108_47# SEL_CONV_TIME[1] 0.00fF
C2471 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C2472 sky130_fd_sc_hd__dfrtn_1_40/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2473 sky130_fd_sc_hd__mux4_2_0/a_1279_413# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C2474 sky130_fd_sc_hd__dfrtn_1_42/a_639_47# RESET_COUNTERn 0.00fF
C2475 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# SEL_CONV_TIME[3] 0.00fF
C2476 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# DOUT[3] 0.30fF
C2477 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__o311a_1_0/a_368_297# 0.00fF
C2478 sky130_fd_sc_hd__inv_1_3/Y DOUT[6] 0.28fF
C2479 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C2480 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_10/a_639_47# 0.00fF
C2481 sky130_fd_sc_hd__inv_1_32/A sky130_fd_sc_hd__inv_1_44/A 0.00fF
C2482 sky130_fd_sc_hd__inv_1_9/Y outb 0.00fF
C2483 sky130_fd_sc_hd__mux4_2_0/a_288_47# sky130_fd_sc_hd__mux4_2_0/a_600_345# -0.00fF
C2484 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtp_1_3/a_651_413# 0.00fF
C2485 sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C2486 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# sky130_fd_sc_hd__dfrtp_1_3/a_543_47# 0.00fF
C2487 sky130_fd_sc_hd__dfrtp_1_2/a_805_47# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C2488 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2489 sky130_fd_sc_hd__nor2_1_0/a_109_297# DOUT[13] 0.00fF
C2490 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# RESET_COUNTERn 0.00fF
C2491 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_2/A 0.02fF
C2492 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C2493 CLK_REF sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C2494 sky130_fd_sc_hd__dfrtn_1_24/a_651_413# SEL_CONV_TIME[0] 0.00fF
C2495 sky130_fd_sc_hd__o221ai_1_0/a_213_123# DOUT[21] 0.00fF
C2496 sky130_fd_sc_hd__nor3_1_14/a_193_297# RESET_COUNTERn 0.00fF
C2497 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__dfrtn_1_34/a_448_47# 0.00fF
C2498 CLK_REF VDD 1.97fF
C2499 sky130_fd_sc_hd__dfrtn_1_31/a_1270_413# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C2500 sky130_fd_sc_hd__dfrtn_1_35/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C2501 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C2502 sky130_fd_sc_hd__inv_1_42/A SEL_CONV_TIME[3] 0.00fF
C2503 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_25/a_193_47# -0.14fF
C2504 DOUT[13] sky130_fd_sc_hd__dfrtn_1_31/a_448_47# 0.01fF
C2505 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_543_47# 0.00fF
C2506 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# 0.00fF
C2507 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__o221ai_1_0/a_295_297# 0.00fF
C2508 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# SEL_CONV_TIME[2] 0.00fF
C2509 SLC_0/a_1235_416# lc_out 0.00fF
C2510 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_29/a_448_47# 0.00fF
C2511 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_1_21/Y 0.14fF
C2512 sky130_fd_sc_hd__nand3b_1_1/a_316_47# SEL_CONV_TIME[3] 0.00fF
C2513 sky130_fd_sc_hd__dfrtn_1_28/a_1283_21# VDD 0.11fF
C2514 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__inv_1_39/Y 0.00fF
C2515 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# -0.00fF
C2516 sky130_fd_sc_hd__dfrtn_1_11/a_761_289# sky130_fd_sc_hd__dfrtn_1_11/a_543_47# -0.00fF
C2517 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# -0.00fF
C2518 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C2519 sky130_fd_sc_hd__or3_1_0/a_183_297# SEL_CONV_TIME[3] 0.00fF
C2520 sky130_fd_sc_hd__dfrtn_1_4/a_761_289# sky130_fd_sc_hd__inv_1_7/Y 0.01fF
C2521 sky130_fd_sc_hd__dfrtn_1_14/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2522 sky130_fd_sc_hd__dfrtn_1_25/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C2523 sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# VDD 0.00fF
C2524 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__inv_1_12/A 0.54fF
C2525 sky130_fd_sc_hd__dfrtn_1_12/a_1217_47# sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# 0.00fF
C2526 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# sky130_fd_sc_hd__dfrtn_1_0/a_1217_47# 0.00fF
C2527 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C2528 sky130_fd_sc_hd__dfrtn_1_16/a_193_47# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C2529 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# DOUT[3] 0.00fF
C2530 sky130_fd_sc_hd__dfrtp_1_0/a_1217_47# RESET_COUNTERn 0.00fF
C2531 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C2532 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__inv_1_37/A 0.01fF
C2533 DOUT[9] sky130_fd_sc_hd__nor3_1_0/a_109_297# 0.00fF
C2534 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# 0.01fF
C2535 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# 0.00fF
C2536 sky130_fd_sc_hd__o221ai_1_0/a_213_123# sky130_fd_sc_hd__o311a_1_0/A3 0.02fF
C2537 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C2538 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.01fF
C2539 DOUT[9] sky130_fd_sc_hd__dfrtn_1_3/a_27_47# 0.00fF
C2540 sky130_fd_sc_hd__dfrtp_1_0/a_639_47# lc_out 0.00fF
C2541 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C2542 sky130_fd_sc_hd__inv_1_2/Y RESET_COUNTERn 0.03fF
C2543 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C2544 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C2545 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C2546 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C2547 sky130_fd_sc_hd__dfrtn_1_39/a_1462_47# RESET_COUNTERn 0.00fF
C2548 sky130_fd_sc_hd__dfrtn_1_20/a_761_289# VDD 0.05fF
C2549 sky130_fd_sc_hd__dfrtn_1_22/a_805_47# sky130_fd_sc_hd__inv_1_39/Y 0.00fF
C2550 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C2551 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C2552 sky130_fd_sc_hd__o311a_1_0/a_266_47# sky130_fd_sc_hd__nand2_1_1/a_113_47# 0.00fF
C2553 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# RESET_COUNTERn -0.03fF
C2554 sky130_fd_sc_hd__dfrtn_1_24/a_448_47# DOUT[21] 0.00fF
C2555 sky130_fd_sc_hd__dfrtn_1_42/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C2556 sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# sky130_fd_sc_hd__inv_1_42/A 0.01fF
C2557 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# DOUT[20] 0.00fF
C2558 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__nor3_1_3/a_109_297# 0.00fF
C2559 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__nand2_1_1/a_113_47# 0.00fF
C2560 sky130_fd_sc_hd__dfrtn_1_18/a_1462_47# RESET_COUNTERn 0.00fF
C2561 sky130_fd_sc_hd__dfrtp_1_3/a_1108_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C2562 DOUT[1] sky130_fd_sc_hd__dfrtn_1_36/a_761_289# 0.00fF
C2563 DOUT[4] sky130_fd_sc_hd__dfrtn_1_8/a_193_47# 0.00fF
C2564 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# SEL_CONV_TIME[0] 0.00fF
C2565 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2566 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_26/a_543_47# 0.01fF
C2567 sky130_fd_sc_hd__dfrtn_1_22/a_1283_21# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C2568 sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2569 sky130_fd_sc_hd__dfrtn_1_42/a_193_47# sky130_fd_sc_hd__dfrtn_1_42/a_761_289# -0.00fF
C2570 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# sky130_fd_sc_hd__dfrtn_1_42/a_543_47# -0.00fF
C2571 sky130_fd_sc_hd__dfrtn_1_30/a_448_47# SEL_CONV_TIME[0] 0.01fF
C2572 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# 0.00fF
C2573 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2574 sky130_fd_sc_hd__mux4_1_0/a_277_47# VDD 0.01fF
C2575 sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C2576 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# DOUT[3] 0.00fF
C2577 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C2578 SLC_0/a_1235_416# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2579 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# VDD 0.01fF
C2580 sky130_fd_sc_hd__dfrtn_1_9/a_639_47# RESET_COUNTERn 0.00fF
C2581 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C2582 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# sky130_fd_sc_hd__dfrtn_1_15/a_761_289# 0.00fF
C2583 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# 0.00fF
C2584 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C2585 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__inv_1_29/Y 0.32fF
C2586 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# DOUT[23] 0.00fF
C2587 sky130_fd_sc_hd__dfrtn_1_24/a_448_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C2588 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C2589 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_193_47# -0.29fF
C2590 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__o221ai_1_0/a_493_297# 0.00fF
C2591 sky130_fd_sc_hd__dfrtn_1_19/a_1270_413# RESET_COUNTERn 0.00fF
C2592 sky130_fd_sc_hd__nor3_1_8/a_109_297# DOUT[7] 0.00fF
C2593 sky130_fd_sc_hd__nor3_1_8/a_193_297# DOUT[6] 0.00fF
C2594 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C2595 sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C2596 CLK_REF sky130_fd_sc_hd__dfrtn_1_17/a_1462_47# 0.00fF
C2597 sky130_fd_sc_hd__nor3_1_4/a_109_297# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C2598 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C2599 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_11/a_27_47# 0.00fF
C2600 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_37/A 0.02fF
C2601 sky130_fd_sc_hd__nor3_1_4/A sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C2602 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C2603 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__inv_1_44/Y 0.01fF
C2604 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# -0.00fF
C2605 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# -0.00fF
C2606 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_6/A 0.02fF
C2607 sky130_fd_sc_hd__dfrtp_1_0/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2608 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# DOUT[20] 0.00fF
C2609 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_4/a_543_47# 0.00fF
C2610 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C2611 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_651_413# 0.00fF
C2612 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C2613 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_4/a_448_47# 0.00fF
C2614 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C2615 sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C2616 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C2617 sky130_fd_sc_hd__dfrtn_1_39/a_193_47# SEL_CONV_TIME[2] 0.00fF
C2618 sky130_fd_sc_hd__nor3_2_3/B DOUT[0] 0.02fF
C2619 sky130_fd_sc_hd__dfrtn_1_11/a_761_289# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C2620 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__inv_1_44/A 0.05fF
C2621 sky130_fd_sc_hd__dfrtn_1_35/a_651_413# sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# 0.00fF
C2622 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# sky130_fd_sc_hd__dfrtn_1_39/a_1462_47# 0.00fF
C2623 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C2624 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C2625 sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C2626 sky130_fd_sc_hd__dfrtn_1_12/a_651_413# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C2627 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_37/a_805_47# 0.00fF
C2628 sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C2629 sky130_fd_sc_hd__dfrtn_1_0/a_1270_413# VDD 0.00fF
C2630 sky130_fd_sc_hd__dfrtn_1_35/a_1283_21# VDD 0.11fF
C2631 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# RESET_COUNTERn 0.05fF
C2632 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__inv_1_15/A 0.05fF
C2633 sky130_fd_sc_hd__inv_1_7/A DOUT[14] 0.02fF
C2634 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# SEL_CONV_TIME[0] 0.01fF
C2635 sky130_fd_sc_hd__dfrtn_1_3/a_1270_413# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C2636 sky130_fd_sc_hd__mux4_2_0/a_27_47# SEL_CONV_TIME[1] -0.00fF
C2637 sky130_fd_sc_hd__inv_1_34/A RESET_COUNTERn 0.62fF
C2638 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# DOUT[19] 0.01fF
C2639 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_38/a_1462_47# 0.00fF
C2640 sky130_fd_sc_hd__dfrtn_1_27/a_543_47# sky130_fd_sc_hd__or3_1_0/C 0.02fF
C2641 SEL_CONV_TIME[0] sky130_fd_sc_hd__inv_1_41/Y 0.04fF
C2642 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# SEL_CONV_TIME[0] 0.00fF
C2643 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_8/Y 0.07fF
C2644 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C2645 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# VDD 0.10fF
C2646 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_14/a_651_413# 0.00fF
C2647 sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C2648 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C2649 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_30/a_761_289# 0.00fF
C2650 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C2651 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__or3b_2_0/B 0.04fF
C2652 sky130_fd_sc_hd__dfrtn_1_39/a_639_47# sky130_fd_sc_hd__inv_1_32/Y 0.00fF
C2653 sky130_fd_sc_hd__inv_1_39/Y RESET_COUNTERn 0.14fF
C2654 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C2655 sky130_fd_sc_hd__or3_1_0/a_111_297# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C2656 sky130_fd_sc_hd__dfrtn_1_24/a_1462_47# RESET_COUNTERn 0.00fF
C2657 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_15/a_543_47# -0.00fF
C2658 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# -0.00fF
C2659 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# -0.00fF
C2660 sky130_fd_sc_hd__dfrtn_1_21/a_639_47# VDD 0.00fF
C2661 sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C2662 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# SLC_0/a_264_22# 0.00fF
C2663 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# SLC_0/a_438_293# 0.00fF
C2664 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# RESET_COUNTERn 0.01fF
C2665 sky130_fd_sc_hd__or3b_2_0/X sky130_fd_sc_hd__o311a_1_0/A3 0.03fF
C2666 sky130_fd_sc_hd__dfrtp_1_0/a_761_289# sky130_fd_sc_hd__inv_1_26/A 0.00fF
C2667 sky130_fd_sc_hd__dfrtn_1_9/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2668 VDD sky130_fd_sc_hd__inv_1_13/A 0.62fF
C2669 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# SEL_CONV_TIME[1] 0.00fF
C2670 sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# sky130_fd_sc_hd__inv_1_40/Y 0.00fF
C2671 CLK_REF sky130_fd_sc_hd__dfrtp_1_3/a_1283_21# 0.01fF
C2672 CLK_REF sky130_fd_sc_hd__o211a_1_0/X 0.00fF
C2673 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_2/a_651_413# 0.00fF
C2674 DOUT[4] sky130_fd_sc_hd__dfrtn_1_8/a_1462_47# 0.00fF
C2675 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# sky130_fd_sc_hd__inv_1_4/Y 0.01fF
C2676 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_4/a_805_47# 0.00fF
C2677 sky130_fd_sc_hd__dfrtn_1_8/a_193_47# outb 0.00fF
C2678 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C2679 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_12/a_651_413# -0.00fF
C2680 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_12/a_448_47# -0.00fF
C2681 sky130_fd_sc_hd__nand3b_1_0/a_232_47# SEL_CONV_TIME[1] 0.00fF
C2682 DOUT[9] sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# 0.00fF
C2683 sky130_fd_sc_hd__dfrtn_1_16/a_805_47# DOUT[2] 0.00fF
C2684 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_651_413# 0.00fF
C2685 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# 0.00fF
C2686 sky130_fd_sc_hd__dfrtn_1_10/a_1283_21# sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# 0.00fF
C2687 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# sky130_fd_sc_hd__dfrtn_1_13/a_193_47# 0.00fF
C2688 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# 0.00fF
C2689 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__dfrtn_1_13/a_761_289# 0.00fF
C2690 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_12/a_193_47# 0.01fF
C2691 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# VIN 0.04fF
C2692 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.01fF
C2693 DOUT[9] sky130_fd_sc_hd__dfrtn_1_4/a_651_413# 0.00fF
C2694 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__inv_1_5/Y 0.01fF
C2695 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# DOUT[11] 0.00fF
C2696 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__dfrtp_1_0/a_448_47# -0.00fF
C2697 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2698 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__inv_1_48/A 0.00fF
C2699 sky130_fd_sc_hd__dfrtn_1_37/a_805_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C2700 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# VIN 0.00fF
C2701 sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C2702 sky130_fd_sc_hd__nor3_1_2/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2703 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__nor3_2_1/a_27_297# 0.00fF
C2704 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C2705 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__nand3b_1_1/Y 0.01fF
C2706 sky130_fd_sc_hd__nor3_1_13/a_109_297# RESET_COUNTERn 0.00fF
C2707 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# DOUT[21] 0.00fF
C2708 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C2709 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# RESET_COUNTERn 0.01fF
C2710 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_11/a_1217_47# 0.00fF
C2711 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# VDD 0.07fF
C2712 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# DOUT[20] 0.00fF
C2713 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# RESET_COUNTERn 0.01fF
C2714 SEL_CONV_TIME[0] sky130_fd_sc_hd__inv_1_49/A 0.04fF
C2715 sky130_fd_sc_hd__dfrtn_1_39/a_1462_47# SEL_CONV_TIME[2] 0.00fF
C2716 sky130_fd_sc_hd__nand3b_1_0/a_53_93# VDD 0.08fF
C2717 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C2718 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# 0.00fF
C2719 sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__inv_1_45/A 0.00fF
C2720 sky130_fd_sc_hd__o311a_1_0/a_81_21# sky130_fd_sc_hd__nor3_1_19/Y -0.00fF
C2721 DOUT[4] sky130_fd_sc_hd__or3b_2_0/B 0.07fF
C2722 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__dfrtn_1_14/a_543_47# 0.00fF
C2723 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_30/a_543_47# 0.00fF
C2724 sky130_fd_sc_hd__dfrtn_1_33/a_448_47# RESET_COUNTERn 0.00fF
C2725 DOUT[1] sky130_fd_sc_hd__dfrtn_1_32/a_639_47# 0.00fF
C2726 sky130_fd_sc_hd__dfrtn_1_7/a_448_47# DOUT[19] 0.00fF
C2727 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__mux4_2_0/a_1060_369# 0.00fF
C2728 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__mux4_2_0/a_1279_413# 0.00fF
C2729 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__mux4_2_0/a_397_47# 0.00fF
C2730 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C2731 sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# RESET_COUNTERn 0.00fF
C2732 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.03fF
C2733 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__inv_1_8/Y 0.01fF
C2734 DOUT[9] sky130_fd_sc_hd__inv_1_14/A 0.00fF
C2735 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# 0.00fF
C2736 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_639_47# 0.00fF
C2737 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__o311a_1_0/A3 0.01fF
C2738 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C2739 sky130_fd_sc_hd__or3_1_0/X sky130_fd_sc_hd__inv_1_42/A 0.00fF
C2740 sky130_fd_sc_hd__mux4_2_0/a_1064_47# SEL_CONV_TIME[1] -0.00fF
C2741 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# DOUT[19] 0.00fF
C2742 DOUT[19] DOUT[8] 0.05fF
C2743 sky130_fd_sc_hd__or3_1_0/a_183_297# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C2744 sky130_fd_sc_hd__dfrtn_1_17/a_543_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C2745 sky130_fd_sc_hd__dfrtp_1_1/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2746 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C2747 sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# VDD 0.00fF
C2748 sky130_fd_sc_hd__nor3_1_16/a_109_297# sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C2749 DOUT[1] sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C2750 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__inv_1_13/A 0.01fF
C2751 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# sky130_fd_sc_hd__inv_1_47/A 0.01fF
C2752 HEADER_0/a_508_138# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C2753 sky130_fd_sc_hd__inv_1_46/Y RESET_COUNTERn 0.02fF
C2754 sky130_fd_sc_hd__dfrtn_1_30/a_639_47# DONE 0.00fF
C2755 sky130_fd_sc_hd__dfrtp_1_0/a_1217_47# SLC_0/a_264_22# 0.00fF
C2756 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C2757 sky130_fd_sc_hd__dfrtn_1_9/a_761_289# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C2758 sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# RESET_COUNTERn 0.03fF
C2759 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.00fF
C2760 sky130_fd_sc_hd__inv_1_6/Y DOUT[14] 0.02fF
C2761 sky130_fd_sc_hd__nand3b_1_0/a_316_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C2762 VDD sky130_fd_sc_hd__inv_1_43/A 0.75fF
C2763 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C2764 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C2765 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.00fF
C2766 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C2767 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.00fF
C2768 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C2769 sky130_fd_sc_hd__dfrtn_1_8/a_1462_47# outb 0.00fF
C2770 sky130_fd_sc_hd__nor3_2_3/a_27_297# RESET_COUNTERn 0.01fF
C2771 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2772 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_10/a_651_413# 0.00fF
C2773 sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C2774 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__inv_1_28/Y 0.09fF
C2775 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_12/a_1462_47# 0.00fF
C2776 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C2777 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__inv_1_27/Y 0.14fF
C2778 sky130_fd_sc_hd__dfrtn_1_24/a_1462_47# SEL_CONV_TIME[3] 0.00fF
C2779 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C2780 sky130_fd_sc_hd__mux4_2_0/a_1060_369# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2781 sky130_fd_sc_hd__mux4_2_0/a_397_47# VDD 0.00fF
C2782 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C2783 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# -0.00fF
C2784 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# -0.00fF
C2785 sky130_fd_sc_hd__dfrtn_1_9/a_761_289# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C2786 sky130_fd_sc_hd__dfrtn_1_21/a_1462_47# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C2787 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# DOUT[14] 0.00fF
C2788 sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# sky130_fd_sc_hd__inv_1_33/A 0.02fF
C2789 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__o311a_1_0/a_266_297# 0.00fF
C2790 sky130_fd_sc_hd__dfrtn_1_27/a_1270_413# SEL_CONV_TIME[1] 0.00fF
C2791 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_2/a_448_47# 0.02fF
C2792 sky130_fd_sc_hd__dfrtn_1_26/a_448_47# RESET_COUNTERn 0.02fF
C2793 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C2794 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__dfrtp_1_3/a_543_47# 0.00fF
C2795 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C2796 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.01fF
C2797 sky130_fd_sc_hd__dfrtn_1_25/a_1270_413# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C2798 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__o211a_1_0/X 0.00fF
C2799 sky130_fd_sc_hd__dfrtn_1_34/a_651_413# RESET_COUNTERn 0.00fF
C2800 sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C2801 sky130_fd_sc_hd__dfrtn_1_35/a_805_47# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C2802 sky130_fd_sc_hd__dfrtn_1_16/a_1108_47# sky130_fd_sc_hd__nor3_2_3/A 0.02fF
C2803 sky130_fd_sc_hd__dfrtn_1_11/a_639_47# VDD 0.00fF
C2804 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2805 sky130_fd_sc_hd__dfrtn_1_19/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# -0.26fF
C2806 sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2807 sky130_fd_sc_hd__dfrtn_1_30/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2808 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C2809 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_37/a_27_47# 0.00fF
C2810 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_37/a_761_289# 0.00fF
C2811 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_37/a_193_47# 0.00fF
C2812 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__inv_1_48/A 0.05fF
C2813 DOUT[2] sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C2814 sky130_fd_sc_hd__dfrtn_1_8/a_651_413# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C2815 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_761_289# 0.00fF
C2816 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C2817 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C2818 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__nor3_2_0/A 0.02fF
C2819 sky130_fd_sc_hd__dfrtn_1_21/a_193_47# sky130_fd_sc_hd__dfrtn_1_19/a_1462_47# 0.00fF
C2820 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_35/a_1283_21# 0.00fF
C2821 sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# DONE 0.00fF
C2822 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.00fF
C2823 sky130_fd_sc_hd__nor3_1_19/Y sky130_fd_sc_hd__or3_1_0/C 0.00fF
C2824 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.01fF
C2825 sky130_fd_sc_hd__mux4_2_0/a_1281_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C2826 sky130_fd_sc_hd__o211a_1_1/a_79_21# DOUT[23] 0.00fF
C2827 sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2828 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C2829 DOUT[9] sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C2830 sky130_fd_sc_hd__dfrtn_1_38/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C2831 sky130_fd_sc_hd__dfrtn_1_27/a_651_413# VDD 0.01fF
C2832 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C2833 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__or2_2_0/a_121_297# 0.00fF
C2834 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_18/a_651_413# 0.00fF
C2835 sky130_fd_sc_hd__nor3_1_18/a_109_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2836 DOUT[1] sky130_fd_sc_hd__dfrtn_1_22/a_27_47# 0.01fF
C2837 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# 0.00fF
C2838 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__dfrtn_1_1/a_448_47# 0.00fF
C2839 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# RESET_COUNTERn 0.00fF
C2840 sky130_fd_sc_hd__nor3_1_19/Y sky130_fd_sc_hd__or2b_1_0/X 0.02fF
C2841 sky130_fd_sc_hd__dfrtn_1_36/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_448_47# -0.00fF
C2842 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_651_413# -0.00fF
C2843 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__nor3_2_0/a_281_297# 0.00fF
C2844 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# DOUT[14] 0.01fF
C2845 sky130_fd_sc_hd__o2111a_2_0/a_458_47# RESET_COUNTERn 0.00fF
C2846 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C2847 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C2848 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C2849 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__a221oi_4_0/a_453_47# -0.00fF
C2850 sky130_fd_sc_hd__dfrtn_1_26/a_651_413# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C2851 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_27_47# 0.00fF
C2852 sky130_fd_sc_hd__dfrtn_1_0/a_543_47# DOUT[18] 0.00fF
C2853 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__inv_1_28/A 0.00fF
C2854 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C2855 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# VDD 0.00fF
C2856 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2857 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.00fF
C2858 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__dfrtn_1_5/a_448_47# 0.00fF
C2859 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C2860 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# sky130_fd_sc_hd__nor3_1_0/A 0.23fF
C2861 VDD DOUT[12] 1.77fF
C2862 sky130_fd_sc_hd__dfrtp_1_3/a_639_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C2863 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C2864 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_27/a_543_47# 0.00fF
C2865 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# SEL_CONV_TIME[1] 0.01fF
C2866 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C2867 sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.03fF
C2868 sky130_fd_sc_hd__dfrtn_1_12/a_805_47# VDD 0.00fF
C2869 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_30/a_1270_413# 0.00fF
C2870 sky130_fd_sc_hd__inv_1_46/Y SEL_CONV_TIME[3] 0.00fF
C2871 sky130_fd_sc_hd__dfrtn_1_14/a_543_47# sky130_fd_sc_hd__nor3_1_1/a_193_297# 0.00fF
C2872 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# sky130_fd_sc_hd__nor3_1_1/a_109_297# 0.00fF
C2873 sky130_fd_sc_hd__dfrtn_1_28/a_1108_47# DOUT[21] 0.00fF
C2874 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# RESET_COUNTERn 0.01fF
C2875 sky130_fd_sc_hd__dfrtn_1_33/a_639_47# DOUT[23] 0.00fF
C2876 sky130_fd_sc_hd__dfrtn_1_39/a_193_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C2877 sky130_fd_sc_hd__dfrtn_1_0/a_1270_413# DOUT[5] 0.00fF
C2878 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__inv_1_50/Y 0.06fF
C2879 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# DOUT[9] 0.00fF
C2880 sky130_fd_sc_hd__dfrtn_1_14/a_651_413# RESET_COUNTERn 0.00fF
C2881 sky130_fd_sc_hd__mux4_1_0/a_757_363# SEL_CONV_TIME[0] 0.01fF
C2882 sky130_fd_sc_hd__dfrtn_1_42/a_639_47# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C2883 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_34/a_805_47# 0.00fF
C2884 sky130_fd_sc_hd__or3b_2_0/a_388_297# SEL_CONV_TIME[1] 0.00fF
C2885 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_42/A 0.02fF
C2886 sky130_fd_sc_hd__inv_1_13/A DOUT[3] 0.00fF
C2887 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# VIN 0.00fF
C2888 sky130_fd_sc_hd__or3_1_0/a_183_297# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C2889 sky130_fd_sc_hd__dfrtn_1_36/a_805_47# sky130_fd_sc_hd__inv_1_40/A 0.00fF
C2890 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C2891 sky130_fd_sc_hd__dfrtn_1_14/a_448_47# DOUT[22] 0.00fF
C2892 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C2893 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C2894 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_13/A 0.16fF
C2895 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# sky130_fd_sc_hd__dfrtn_1_37/a_543_47# 0.00fF
C2896 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__dfrtn_1_37/a_1270_413# 0.00fF
C2897 sky130_fd_sc_hd__dfrtn_1_40/a_1270_413# sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# 0.00fF
C2898 sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# sky130_fd_sc_hd__dfrtn_1_37/a_761_289# 0.00fF
C2899 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_37/a_448_47# 0.00fF
C2900 sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C2901 DOUT[1] sky130_fd_sc_hd__dfrtn_1_23/a_193_47# 0.00fF
C2902 sky130_fd_sc_hd__dfrtn_1_40/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2903 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__inv_1_27/Y 0.01fF
C2904 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__nor3_2_3/C -0.03fF
C2905 sky130_fd_sc_hd__a221oi_4_0/a_453_47# VDD 0.01fF
C2906 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# 0.00fF
C2907 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C2908 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# 0.00fF
C2909 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C2910 sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# SEL_CONV_TIME[2] 0.00fF
C2911 sky130_fd_sc_hd__dfrtn_1_22/a_1108_47# sky130_fd_sc_hd__inv_1_39/A 0.01fF
C2912 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_24/a_639_47# -0.00fF
C2913 sky130_fd_sc_hd__mux4_1_0/X RESET_COUNTERn 0.01fF
C2914 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2915 sky130_fd_sc_hd__dfrtn_1_42/a_651_413# DOUT[2] 0.00fF
C2916 VDD sky130_fd_sc_hd__inv_1_3/A 0.58fF
C2917 sky130_fd_sc_hd__o221ai_1_0/a_295_297# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C2918 sky130_fd_sc_hd__nor3_1_12/a_109_297# VDD 0.00fF
C2919 sky130_fd_sc_hd__or3b_2_0/a_27_47# VDD 0.06fF
C2920 sky130_fd_sc_hd__dfrtn_1_39/a_639_47# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C2921 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# -0.00fF
C2922 DOUT[1] sky130_fd_sc_hd__dfrtn_1_22/a_1217_47# 0.00fF
C2923 sky130_fd_sc_hd__dfrtn_1_31/a_761_289# SEL_CONV_TIME[1] 0.00fF
C2924 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C2925 DOUT[4] sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C2926 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# RESET_COUNTERn 0.00fF
C2927 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_41/a_651_413# 0.00fF
C2928 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_19/a_1283_21# 0.02fF
C2929 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_31/a_27_47# 0.00fF
C2930 sky130_fd_sc_hd__dfrtn_1_26/a_639_47# DOUT[23] 0.00fF
C2931 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# DOUT[19] 0.01fF
C2932 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# DOUT[14] 0.00fF
C2933 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_15/a_651_413# 0.00fF
C2934 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_805_47# 0.00fF
C2935 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_639_47# 0.00fF
C2936 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C2937 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# 0.00fF
C2938 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__dfrtn_1_15/a_543_47# 0.00fF
C2939 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# 0.00fF
C2940 sky130_fd_sc_hd__dfrtn_1_5/a_805_47# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C2941 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# 0.00fF
C2942 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C2943 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C2944 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_639_47# 0.00fF
C2945 sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C2946 sky130_fd_sc_hd__dfrtn_1_17/a_543_47# VDD 0.05fF
C2947 sky130_fd_sc_hd__dfrtn_1_17/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2948 sky130_fd_sc_hd__inv_1_36/A sky130_fd_sc_hd__inv_1_40/Y 0.00fF
C2949 sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# sky130_fd_sc_hd__inv_1_8/A 0.01fF
C2950 sky130_fd_sc_hd__dfrtn_1_36/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C2951 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C2952 sky130_fd_sc_hd__dfrtn_1_36/a_805_47# VDD 0.00fF
C2953 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# 0.00fF
C2954 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# 0.00fF
C2955 sky130_fd_sc_hd__dfrtn_1_12/a_651_413# sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# 0.00fF
C2956 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__o2111a_2_0/a_674_297# 0.00fF
C2957 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__o2111a_2_0/a_80_21# 0.00fF
C2958 sky130_fd_sc_hd__or3_1_0/a_111_297# sky130_fd_sc_hd__o2111a_2_0/a_80_21# 0.00fF
C2959 sky130_fd_sc_hd__dfrtn_1_21/a_193_47# sky130_fd_sc_hd__dfrtn_1_21/a_543_47# -0.00fF
C2960 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# 0.00fF
C2961 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C2962 sky130_fd_sc_hd__dfrtn_1_0/a_1462_47# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C2963 sky130_fd_sc_hd__dfrtn_1_17/a_805_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C2964 DOUT[9] VIN 0.01fF
C2965 VDD sky130_fd_sc_hd__nor3_2_3/C 11.78fF
C2966 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C2967 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C2968 sky130_fd_sc_hd__o2111a_2_0/a_458_47# SEL_CONV_TIME[3] 0.00fF
C2969 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C2970 sky130_fd_sc_hd__o311a_1_0/a_368_297# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C2971 sky130_fd_sc_hd__o211a_1_0/a_79_21# DOUT[15] 0.02fF
C2972 sky130_fd_sc_hd__dfrtp_1_0/a_1283_21# outb 0.00fF
C2973 sky130_fd_sc_hd__o311a_1_0/a_81_21# SEL_CONV_TIME[0] 0.00fF
C2974 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__nand3b_1_1/a_53_93# 0.00fF
C2975 sky130_fd_sc_hd__dfrtn_1_28/a_1217_47# RESET_COUNTERn 0.00fF
C2976 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# VDD 0.11fF
C2977 sky130_fd_sc_hd__dfrtn_1_39/a_1462_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C2978 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__nor3_1_1/a_193_297# 0.00fF
C2979 sky130_fd_sc_hd__mux4_2_0/a_372_413# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C2980 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# sky130_fd_sc_hd__nor3_1_1/a_109_297# 0.00fF
C2981 sky130_fd_sc_hd__mux4_2_0/a_193_369# SEL_CONV_TIME[0] 0.00fF
C2982 sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# RESET_COUNTERn 0.03fF
C2983 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# RESET_COUNTERn 0.02fF
C2984 sky130_fd_sc_hd__dfrtn_1_35/a_1108_47# DOUT[21] 0.00fF
C2985 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_12/a_448_47# 0.00fF
C2986 sky130_fd_sc_hd__dfrtn_1_3/a_1270_413# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C2987 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C2988 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__inv_1_1/Y 0.16fF
C2989 sky130_fd_sc_hd__dfrtn_1_23/a_448_47# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C2990 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C2991 sky130_fd_sc_hd__dfrtn_1_18/a_1462_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C2992 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# 0.00fF
C2993 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_39/a_193_47# 0.00fF
C2994 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_651_413# 0.00fF
C2995 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# 0.00fF
C2996 sky130_fd_sc_hd__nor3_1_4/a_193_297# VDD 0.00fF
C2997 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__inv_1_33/A 0.00fF
C2998 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C2999 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# 0.00fF
C3000 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C3001 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_19/a_543_47# 0.00fF
C3002 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C3003 DOUT[13] sky130_fd_sc_hd__nand2_1_2/Y 0.00fF
C3004 sky130_fd_sc_hd__inv_1_45/Y SEL_CONV_TIME[0] 0.01fF
C3005 sky130_fd_sc_hd__dfrtn_1_32/a_805_47# sky130_fd_sc_hd__inv_1_9/A 0.00fF
C3006 sky130_fd_sc_hd__dfrtn_1_0/a_543_47# DOUT[22] 0.00fF
C3007 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__inv_1_31/A 0.01fF
C3008 sky130_fd_sc_hd__dfrtn_1_21/a_193_47# sky130_fd_sc_hd__inv_1_35/Y 0.11fF
C3009 sky130_fd_sc_hd__dfrtn_1_20/a_639_47# RESET_COUNTERn 0.00fF
C3010 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# SEL_CONV_TIME[0] 0.00fF
C3011 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C3012 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__o221ai_1_0/a_295_297# 0.00fF
C3013 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__o221ai_1_0/a_493_297# 0.00fF
C3014 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_38/a_543_47# 0.00fF
C3015 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__inv_1_29/Y 0.00fF
C3016 DOUT[1] sky130_fd_sc_hd__dfrtn_1_23/a_1462_47# 0.00fF
C3017 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.00fF
C3018 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C3019 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_651_413# 0.00fF
C3020 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# 0.00fF
C3021 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C3022 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_448_47# 0.00fF
C3023 sky130_fd_sc_hd__dfrtn_1_18/a_805_47# DOUT[2] 0.00fF
C3024 sky130_fd_sc_hd__o2111a_2_0/a_458_47# SEL_CONV_TIME[2] 0.00fF
C3025 sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# sky130_fd_sc_hd__inv_1_25/A 0.00fF
C3026 sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3027 sky130_fd_sc_hd__dfrtn_1_32/a_448_47# VDD 0.01fF
C3028 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C3029 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# sky130_fd_sc_hd__inv_1_6/Y 0.10fF
C3030 DOUT[11] sky130_fd_sc_hd__nor3_2_3/B 0.07fF
C3031 sky130_fd_sc_hd__nor3_2_1/a_281_297# VDD 0.04fF
C3032 DOUT[23] sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C3033 sky130_fd_sc_hd__nand3b_1_0/a_316_47# SEL_CONV_TIME[0] 0.00fF
C3034 sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C3035 sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C3036 sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# sky130_fd_sc_hd__inv_1_52/Y 0.02fF
C3037 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C3038 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_1462_47# 0.00fF
C3039 sky130_fd_sc_hd__dfrtp_1_3/a_761_289# sky130_fd_sc_hd__or2_2_0/A 0.02fF
C3040 sky130_fd_sc_hd__inv_1_36/A sky130_fd_sc_hd__inv_1_36/Y 0.01fF
C3041 sky130_fd_sc_hd__mux4_2_0/a_27_47# DOUT[21] 0.00fF
C3042 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# 0.00fF
C3043 sky130_fd_sc_hd__mux4_1_0/a_193_47# RESET_COUNTERn 0.00fF
C3044 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__inv_1_37/A 0.01fF
C3045 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C3046 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__inv_1_2/Y 0.01fF
C3047 sky130_fd_sc_hd__inv_1_12/A sky130_fd_sc_hd__inv_1_8/Y 0.02fF
C3048 sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# sky130_fd_sc_hd__dfrtn_1_28/a_27_47# 0.02fF
C3049 sky130_fd_sc_hd__o211a_1_0/a_510_47# RESET_COUNTERn 0.00fF
C3050 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# 0.00fF
C3051 sky130_fd_sc_hd__mux4_1_0/X SEL_CONV_TIME[3] 0.28fF
C3052 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C3053 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_805_47# 0.00fF
C3054 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_31/a_1217_47# 0.00fF
C3055 sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# sky130_fd_sc_hd__o2111a_2_0/X 0.01fF
C3056 sky130_fd_sc_hd__dfrtn_1_34/a_448_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C3057 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C3058 sky130_fd_sc_hd__o211a_1_0/a_297_297# lc_out 0.00fF
C3059 sky130_fd_sc_hd__dfrtn_1_28/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3060 sky130_fd_sc_hd__dfrtn_1_42/a_761_289# sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C3061 sky130_fd_sc_hd__inv_1_10/A DOUT[12] 0.00fF
C3062 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# DOUT[11] 0.00fF
C3063 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# DOUT[9] 0.00fF
C3064 sky130_fd_sc_hd__dfrtn_1_32/a_193_47# sky130_fd_sc_hd__dfrtn_1_32/a_639_47# -0.00fF
C3065 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# VDD 0.05fF
C3066 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C3067 sky130_fd_sc_hd__dfrtn_1_0/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3068 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__inv_1_33/A 0.01fF
C3069 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_34/a_27_47# 0.00fF
C3070 sky130_fd_sc_hd__dfrtn_1_22/a_805_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C3071 sky130_fd_sc_hd__inv_1_15/A sky130_fd_sc_hd__nor3_1_0/A 0.04fF
C3072 DOUT[4] sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# 0.00fF
C3073 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__dfrtn_1_30/a_651_413# -0.00fF
C3074 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__dfrtn_1_30/a_448_47# -0.00fF
C3075 sky130_fd_sc_hd__nand3b_1_0/a_232_47# DOUT[21] 0.00fF
C3076 sky130_fd_sc_hd__nor3_1_9/a_193_297# DOUT[11] 0.00fF
C3077 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C3078 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_805_47# 0.00fF
C3079 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C3080 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_639_47# 0.00fF
C3081 sky130_fd_sc_hd__nor3_1_5/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3082 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C3083 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C3084 sky130_fd_sc_hd__nor3_1_11/a_193_297# sky130_fd_sc_hd__dfrtn_1_7/a_448_47# 0.00fF
C3085 sky130_fd_sc_hd__dfrtn_1_19/a_193_47# sky130_fd_sc_hd__inv_1_28/A 0.46fF
C3086 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfrtn_1_41/a_651_413# 0.00fF
C3087 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__inv_1_8/Y 0.05fF
C3088 sky130_fd_sc_hd__dfrtn_1_31/a_1462_47# VDD 0.00fF
C3089 sky130_fd_sc_hd__inv_1_52/A DOUT[13] 0.01fF
C3090 sky130_fd_sc_hd__dfrtn_1_3/a_651_413# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C3091 sky130_fd_sc_hd__mux4_1_0/X SEL_CONV_TIME[2] 0.00fF
C3092 SEL_CONV_TIME[0] sky130_fd_sc_hd__or3_1_0/C 0.02fF
C3093 sky130_fd_sc_hd__dfrtn_1_28/a_651_413# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C3094 sky130_fd_sc_hd__mux4_2_0/a_1281_47# SEL_CONV_TIME[0] 0.00fF
C3095 sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C3096 sky130_fd_sc_hd__dfrtn_1_32/a_27_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C3097 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C3098 sky130_fd_sc_hd__dfrtn_1_35/a_1217_47# RESET_COUNTERn -0.00fF
C3099 DOUT[9] sky130_fd_sc_hd__inv_1_1/A 0.00fF
C3100 sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C3101 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_1217_47# -0.00fF
C3102 CLK_REF sky130_fd_sc_hd__dfrtn_1_21/a_193_47# 0.02fF
C3103 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_1/a_27_47# 0.00fF
C3104 sky130_fd_sc_hd__nor3_1_11/a_109_297# RESET_COUNTERn 0.00fF
C3105 sky130_fd_sc_hd__nor3_1_11/a_193_297# DOUT[8] 0.00fF
C3106 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_8/A 0.01fF
C3107 sky130_fd_sc_hd__or2b_1_0/X SEL_CONV_TIME[0] 0.96fF
C3108 sky130_fd_sc_hd__nand3b_1_1/Y sky130_fd_sc_hd__inv_1_44/Y 0.10fF
C3109 sky130_fd_sc_hd__nor3_1_8/a_109_297# VIN 0.00fF
C3110 sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# RESET_COUNTERn 0.00fF
C3111 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_25/a_27_47# 0.00fF
C3112 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__dfrtn_1_25/a_193_47# 0.00fF
C3113 sky130_fd_sc_hd__dfrtp_1_3/a_761_289# sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# 0.00fF
C3114 sky130_fd_sc_hd__dfrtp_1_3/a_543_47# sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# 0.00fF
C3115 sky130_fd_sc_hd__dfrtp_1_3/a_448_47# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C3116 sky130_fd_sc_hd__dfrtn_1_4/a_805_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C3117 sky130_fd_sc_hd__o2111a_2_0/a_386_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C3118 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C3119 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__inv_1_43/Y 0.01fF
C3120 sky130_fd_sc_hd__dfrtn_1_34/a_639_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C3121 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C3122 sky130_fd_sc_hd__nand3b_1_0/a_232_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C3123 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_18/a_1462_47# 0.00fF
C3124 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C3125 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_7/A 0.02fF
C3126 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__dfrtn_1_29/a_448_47# 0.00fF
C3127 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# 0.00fF
C3128 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__dfrtn_1_29/a_651_413# 0.00fF
C3129 sky130_fd_sc_hd__dfrtn_1_4/a_543_47# sky130_fd_sc_hd__inv_1_7/A 0.01fF
C3130 sky130_fd_sc_hd__dfrtn_1_10/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3131 sky130_fd_sc_hd__o211a_1_0/a_297_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3132 sky130_fd_sc_hd__nand2_1_0/a_113_47# outb 0.00fF
C3133 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C3134 sky130_fd_sc_hd__dfrtp_1_3/a_448_47# VDD 0.01fF
C3135 sky130_fd_sc_hd__dfrtp_1_3/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3136 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__o211a_1_0/X 0.15fF
C3137 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__nor3_1_12/a_109_297# 0.00fF
C3138 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_1/a_639_47# -0.00fF
C3139 sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# SEL_CONV_TIME[1] 0.00fF
C3140 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C3141 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C3142 sky130_fd_sc_hd__or3b_2_0/a_388_297# sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# 0.00fF
C3143 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# 0.00fF
C3144 DOUT[4] sky130_fd_sc_hd__dfrtn_1_34/a_27_47# 0.02fF
C3145 sky130_fd_sc_hd__mux4_2_0/a_193_47# RESET_COUNTERn 0.00fF
C3146 sky130_fd_sc_hd__dfrtn_1_23/a_1217_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C3147 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__dfrtp_1_1/D 0.00fF
C3148 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.06fF
C3149 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_36/a_805_47# 0.00fF
C3150 sky130_fd_sc_hd__inv_1_44/Y sky130_fd_sc_hd__inv_1_51/Y 0.01fF
C3151 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_543_47# -0.00fF
C3152 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# -0.00fF
C3153 sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# RESET_COUNTERn 0.01fF
C3154 sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# DOUT[11] 0.00fF
C3155 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__nor3_2_3/C 0.37fF
C3156 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_10/a_27_47# 0.01fF
C3157 sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# DOUT[9] 0.00fF
C3158 sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3159 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# DOUT[23] 0.00fF
C3160 sky130_fd_sc_hd__dfrtn_1_35/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3161 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# DOUT[19] 0.00fF
C3162 sky130_fd_sc_hd__nor3_1_15/a_193_297# VDD 0.00fF
C3163 sky130_fd_sc_hd__dfrtn_1_8/a_27_47# DOUT[12] 0.02fF
C3164 sky130_fd_sc_hd__dfrtn_1_41/a_805_47# RESET_COUNTERn 0.00fF
C3165 sky130_fd_sc_hd__inv_1_3/A DOUT[3] 0.00fF
C3166 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_34/a_1217_47# 0.00fF
C3167 sky130_fd_sc_hd__inv_1_37/A RESET_COUNTERn 0.40fF
C3168 sky130_fd_sc_hd__dfrtn_1_18/a_27_47# sky130_fd_sc_hd__inv_1_27/Y 0.00fF
C3169 sky130_fd_sc_hd__nor3_2_1/a_281_297# sky130_fd_sc_hd__o211a_1_0/X 0.00fF
C3170 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C3171 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# VDD 0.01fF
C3172 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__o2111a_2_0/X 0.01fF
C3173 sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C3174 sky130_fd_sc_hd__dfrtp_1_1/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3175 CLK_REF sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.02fF
C3176 sky130_fd_sc_hd__nor3_2_3/a_27_297# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C3177 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_3/A 0.04fF
C3178 sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C3179 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.00fF
C3180 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__inv_1_47/Y 0.00fF
C3181 sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.00fF
C3182 sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# sky130_fd_sc_hd__dfrtn_1_18/a_761_289# 0.01fF
C3183 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_448_47# 0.00fF
C3184 CLK_REF sky130_fd_sc_hd__inv_1_29/Y 0.00fF
C3185 sky130_fd_sc_hd__dfrtn_1_32/a_1217_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C3186 sky130_fd_sc_hd__nor3_1_1/a_109_297# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C3187 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_34/a_27_47# 0.00fF
C3188 sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C3189 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_448_47# 0.00fF
C3190 sky130_fd_sc_hd__dfrtn_1_23/a_543_47# sky130_fd_sc_hd__dfrtn_1_36/a_543_47# 0.00fF
C3191 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# sky130_fd_sc_hd__dfrtn_1_36/a_761_289# 0.00fF
C3192 sky130_fd_sc_hd__dfrtn_1_27/a_543_47# RESET_COUNTERn 0.01fF
C3193 sky130_fd_sc_hd__dfrtn_1_27/a_1270_413# DOUT[21] 0.00fF
C3194 sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C3195 sky130_fd_sc_hd__o2111a_2_0/a_458_47# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C3196 sky130_fd_sc_hd__dfrtn_1_35/a_1283_21# sky130_fd_sc_hd__inv_1_38/A 0.01fF
C3197 sky130_fd_sc_hd__dfrtn_1_3/a_639_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C3198 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C3199 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__inv_1_49/A 0.02fF
C3200 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__dfrtn_1_25/a_448_47# 0.00fF
C3201 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__dfrtn_1_25/a_651_413# 0.00fF
C3202 sky130_fd_sc_hd__dfrtp_1_3/a_651_413# sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# 0.00fF
C3203 sky130_fd_sc_hd__nor3_2_3/C DOUT[3] 0.19fF
C3204 sky130_fd_sc_hd__nor3_2_0/a_27_297# sky130_fd_sc_hd__dfrtn_1_12/a_193_47# 0.00fF
C3205 sky130_fd_sc_hd__nor3_2_0/a_281_297# sky130_fd_sc_hd__dfrtn_1_12/a_27_47# 0.00fF
C3206 sky130_fd_sc_hd__o311a_1_0/a_266_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3207 sky130_fd_sc_hd__dfrtn_1_38/a_761_289# DOUT[2] 0.00fF
C3208 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C3209 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# sky130_fd_sc_hd__mux4_2_0/a_600_345# 0.00fF
C3210 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# sky130_fd_sc_hd__mux4_2_0/a_872_316# 0.00fF
C3211 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.00fF
C3212 sky130_fd_sc_hd__dfrtn_1_37/a_639_47# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C3213 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# sky130_fd_sc_hd__mux4_2_0/a_193_47# 0.00fF
C3214 sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C3215 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C3216 sky130_fd_sc_hd__dfrtn_1_4/a_651_413# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C3217 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3218 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C3219 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# sky130_fd_sc_hd__nor3_1_2/a_193_297# 0.00fF
C3220 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C3221 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# DOUT[21] 0.02fF
C3222 sky130_fd_sc_hd__dfrtn_1_29/a_639_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C3223 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__inv_1_32/A 0.84fF
C3224 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__nor3_2_3/C 0.17fF
C3225 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# RESET_COUNTERn 0.02fF
C3226 sky130_fd_sc_hd__dfrtn_1_9/a_761_289# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C3227 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__or3_1_0/X 0.01fF
C3228 sky130_fd_sc_hd__dfrtn_1_33/a_543_47# sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# 0.00fF
C3229 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# 0.00fF
C3230 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__inv_1_0/Y 0.02fF
C3231 DOUT[5] sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C3232 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C3233 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# VDD 0.18fF
C3234 sky130_fd_sc_hd__dfrtn_1_22/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3235 sky130_fd_sc_hd__dfrtn_1_39/a_761_289# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C3236 sky130_fd_sc_hd__dfrtn_1_22/a_1270_413# VDD 0.00fF
C3237 DOUT[1] sky130_fd_sc_hd__dfrtn_1_42/a_448_47# 0.00fF
C3238 sky130_fd_sc_hd__nor3_1_12/a_109_297# sky130_fd_sc_hd__dfrtn_1_8/a_27_47# 0.00fF
C3239 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3240 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# RESET_COUNTERn 0.01fF
C3241 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# -0.00fF
C3242 sky130_fd_sc_hd__dfrtn_1_38/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_543_47# -0.00fF
C3243 sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C3244 sky130_fd_sc_hd__nor3_1_5/A RESET_COUNTERn 0.29fF
C3245 sky130_fd_sc_hd__dfrtn_1_28/a_805_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C3246 sky130_fd_sc_hd__nor3_1_20/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3247 sky130_fd_sc_hd__dfrtn_1_41/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3248 sky130_fd_sc_hd__nor3_1_4/a_193_297# DOUT[3] 0.00fF
C3249 DOUT[4] sky130_fd_sc_hd__dfrtn_1_34/a_1217_47# 0.00fF
C3250 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__dfrtn_1_25/a_27_47# 0.00fF
C3251 sky130_fd_sc_hd__or3b_2_0/a_472_297# SEL_CONV_TIME[0] 0.00fF
C3252 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C3253 sky130_fd_sc_hd__dfrtn_1_18/a_761_289# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C3254 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_1_17/A 0.04fF
C3255 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C3256 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__inv_1_28/A 0.00fF
C3257 sky130_fd_sc_hd__dfrtn_1_23/a_639_47# sky130_fd_sc_hd__inv_1_40/A 0.00fF
C3258 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# 0.00fF
C3259 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# sky130_fd_sc_hd__dfrtp_1_1/a_193_47# 0.00fF
C3260 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/a_543_47# 0.00fF
C3261 sky130_fd_sc_hd__nor3_1_4/a_193_297# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C3262 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C3263 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.00fF
C3264 sky130_fd_sc_hd__o211a_1_1/a_297_297# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C3265 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_26/a_761_289# 0.00fF
C3266 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__inv_1_42/Y 0.01fF
C3267 sky130_fd_sc_hd__dfrtn_1_8/a_448_47# sky130_fd_sc_hd__inv_1_9/A 0.00fF
C3268 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_10/a_1217_47# 0.00fF
C3269 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C3270 sky130_fd_sc_hd__dfrtn_1_26/a_761_289# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C3271 sky130_fd_sc_hd__dfrtn_1_26/a_448_47# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C3272 sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# DOUT[23] 0.00fF
C3273 sky130_fd_sc_hd__dfrtn_1_8/a_1217_47# DOUT[12] 0.00fF
C3274 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# sky130_fd_sc_hd__inv_1_5/A 0.02fF
C3275 sky130_fd_sc_hd__dfrtn_1_3/a_1270_413# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C3276 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C3277 sky130_fd_sc_hd__mux4_2_0/a_193_47# SEL_CONV_TIME[3] 0.00fF
C3278 sky130_fd_sc_hd__nor3_2_1/A SLC_0/a_919_243# 0.00fF
C3279 sky130_fd_sc_hd__dfrtn_1_27/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.03fF
C3280 sky130_fd_sc_hd__dfrtn_1_16/a_448_47# VDD 0.01fF
C3281 sky130_fd_sc_hd__dfrtn_1_16/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.04fF
C3282 sky130_fd_sc_hd__or3_1_0/X sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C3283 SLC_0/a_264_22# sky130_fd_sc_hd__o211a_1_0/a_510_47# 0.00fF
C3284 sky130_fd_sc_hd__dfrtn_1_8/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.04fF
C3285 sky130_fd_sc_hd__dfrtn_1_8/a_761_289# VDD 0.05fF
C3286 sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C3287 sky130_fd_sc_hd__dfrtn_1_18/a_1217_47# sky130_fd_sc_hd__inv_1_27/Y 0.00fF
C3288 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# -0.28fF
C3289 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C3290 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_639_47# -0.00fF
C3291 sky130_fd_sc_hd__inv_1_14/A sky130_fd_sc_hd__inv_1_8/Y 0.01fF
C3292 sky130_fd_sc_hd__dfrtn_1_7/a_543_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C3293 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# DOUT[21] 0.00fF
C3294 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__inv_1_47/A 0.01fF
C3295 CLK_REF sky130_fd_sc_hd__dfrtn_1_19/a_1217_47# 0.00fF
C3296 sky130_fd_sc_hd__dfrtn_1_21/a_651_413# sky130_fd_sc_hd__inv_1_35/A 0.00fF
C3297 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# 0.02fF
C3298 sky130_fd_sc_hd__dfrtn_1_20/a_1217_47# sky130_fd_sc_hd__dfrtn_1_18/a_448_47# 0.00fF
C3299 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C3300 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__dfrtn_1_29/a_805_47# 0.00fF
C3301 sky130_fd_sc_hd__dfrtn_1_18/a_805_47# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C3302 sky130_fd_sc_hd__dfrtn_1_31/a_543_47# SEL_CONV_TIME[0] 0.01fF
C3303 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C3304 sky130_fd_sc_hd__dfrtp_1_0/a_1270_413# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C3305 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C3306 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# -0.00fF
C3307 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# -0.00fF
C3308 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_40/a_543_47# -0.00fF
C3309 sky130_fd_sc_hd__inv_1_3/A DOUT[20] 0.00fF
C3310 sky130_fd_sc_hd__nor3_2_1/A out 0.01fF
C3311 sky130_fd_sc_hd__dfrtn_1_23/a_1217_47# sky130_fd_sc_hd__dfrtn_1_36/a_448_47# 0.00fF
C3312 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C3313 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__inv_1_13/A 0.00fF
C3314 sky130_fd_sc_hd__o211a_1_0/a_215_47# out 0.00fF
C3315 sky130_fd_sc_hd__nor3_1_12/a_193_297# DOUT[21] 0.00fF
C3316 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__inv_1_13/Y 0.01fF
C3317 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3318 sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# sky130_fd_sc_hd__nor3_2_0/A 0.01fF
C3319 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__inv_1_44/A 0.00fF
C3320 sky130_fd_sc_hd__dfrtn_1_9/a_543_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C3321 sky130_fd_sc_hd__mux4_2_0/a_193_47# SEL_CONV_TIME[2] 0.00fF
C3322 sky130_fd_sc_hd__nor3_1_11/a_109_297# sky130_fd_sc_hd__dfrtn_1_2/a_448_47# 0.00fF
C3323 sky130_fd_sc_hd__dfrtn_1_9/a_805_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C3324 sky130_fd_sc_hd__dfrtn_1_23/a_639_47# VDD 0.00fF
C3325 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3326 sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C3327 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_35/a_1270_413# 0.00fF
C3328 DOUT[13] sky130_fd_sc_hd__dfrtn_1_30/a_805_47# 0.00fF
C3329 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_639_47# 0.00fF
C3330 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_805_47# 0.00fF
C3331 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C3332 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C3333 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__o311a_1_0/A3 0.03fF
C3334 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_3/a_761_289# 0.00fF
C3335 sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# VDD 0.05fF
C3336 sky130_fd_sc_hd__dfrtn_1_7/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3337 sky130_fd_sc_hd__inv_1_45/A SEL_CONV_TIME[0] 0.12fF
C3338 sky130_fd_sc_hd__dfrtn_1_42/a_1217_47# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C3339 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# DOUT[14] 0.01fF
C3340 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__inv_1_29/Y 0.00fF
C3341 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C3342 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_13/A 0.00fF
C3343 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__inv_1_5/Y 0.10fF
C3344 sky130_fd_sc_hd__dfrtn_1_36/a_448_47# RESET_COUNTERn 0.01fF
C3345 sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# DOUT[21] 0.00fF
C3346 sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C3347 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C3348 DOUT[4] sky130_fd_sc_hd__dfrtn_1_28/a_1283_21# 0.01fF
C3349 sky130_fd_sc_hd__dfrtp_1_0/a_1270_413# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C3350 sky130_fd_sc_hd__or2_2_0/B out 0.00fF
C3351 sky130_fd_sc_hd__o311a_1_0/a_266_47# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C3352 sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C3353 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3354 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# VDD 0.00fF
C3355 VDD DOUT[7] 0.93fF
C3356 sky130_fd_sc_hd__nor3_2_3/C DOUT[20] 0.07fF
C3357 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C3358 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C3359 sky130_fd_sc_hd__or3b_2_0/a_388_297# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C3360 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C3361 sky130_fd_sc_hd__or2b_1_0/a_219_297# SEL_CONV_TIME[0] 0.04fF
C3362 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C3363 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C3364 sky130_fd_sc_hd__inv_1_50/A VDD 0.47fF
C3365 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C3366 sky130_fd_sc_hd__dfrtn_1_27/a_448_47# DOUT[23] 0.00fF
C3367 sky130_fd_sc_hd__dfrtp_1_0/a_805_47# sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# 0.00fF
C3368 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# 0.00fF
C3369 sky130_fd_sc_hd__dfrtp_1_1/a_448_47# DOUT[0] 0.00fF
C3370 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C3371 sky130_fd_sc_hd__nor3_1_18/a_193_297# DOUT[23] 0.00fF
C3372 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C3373 CLK_REF sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.03fF
C3374 sky130_fd_sc_hd__inv_1_33/A sky130_fd_sc_hd__inv_1_44/A 0.01fF
C3375 sky130_fd_sc_hd__inv_1_53/A sky130_fd_sc_hd__mux4_1_0/X 0.01fF
C3376 sky130_fd_sc_hd__inv_1_43/Y SEL_CONV_TIME[1] 0.01fF
C3377 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# SEL_CONV_TIME[1] 0.00fF
C3378 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_651_413# 0.00fF
C3379 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# 0.00fF
C3380 sky130_fd_sc_hd__dfrtn_1_25/a_651_413# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C3381 sky130_fd_sc_hd__dfrtn_1_25/a_448_47# sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.00fF
C3382 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# 0.00fF
C3383 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_15/A 0.00fF
C3384 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C3385 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C3386 sky130_fd_sc_hd__dfrtn_1_26/a_448_47# sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# 0.00fF
C3387 sky130_fd_sc_hd__dfrtn_1_42/a_1108_47# sky130_fd_sc_hd__inv_1_37/A 0.01fF
C3388 sky130_fd_sc_hd__nor3_1_4/a_193_297# DOUT[20] 0.00fF
C3389 sky130_fd_sc_hd__nor3_1_4/a_109_297# DOUT[6] 0.00fF
C3390 DOUT[9] sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C3391 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C3392 sky130_fd_sc_hd__dfrtn_1_27/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3393 sky130_fd_sc_hd__dfrtn_1_8/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3394 sky130_fd_sc_hd__nor3_1_14/a_109_297# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C3395 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C3396 DOUT[9] DOUT[17] 0.10fF
C3397 sky130_fd_sc_hd__dfrtn_1_34/a_1270_413# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C3398 VDD sky130_fd_sc_hd__inv_1_12/A 0.73fF
C3399 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C3400 sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C3401 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C3402 sky130_fd_sc_hd__dfrtn_1_23/a_543_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C3403 sky130_fd_sc_hd__dfrtn_1_32/a_761_289# RESET_COUNTERn 0.00fF
C3404 sky130_fd_sc_hd__nor3_1_19/Y RESET_COUNTERn 0.02fF
C3405 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__dfrtn_1_33/a_27_47# 0.00fF
C3406 sky130_fd_sc_hd__dfrtn_1_8/a_193_47# sky130_fd_sc_hd__inv_1_9/Y 0.18fF
C3407 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__inv_1_42/Y 0.01fF
C3408 sky130_fd_sc_hd__dfrtp_1_2/a_448_47# CLK_REF 0.00fF
C3409 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__or3b_2_0/a_176_21# 0.03fF
C3410 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__dfrtn_1_22/a_543_47# -0.00fF
C3411 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# sky130_fd_sc_hd__dfrtn_1_22/a_761_289# -0.00fF
C3412 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_21/a_27_47# 0.00fF
C3413 sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3414 sky130_fd_sc_hd__or2b_1_0/a_301_297# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C3415 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C3416 sky130_fd_sc_hd__inv_1_9/A sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3417 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# sky130_fd_sc_hd__inv_1_44/A 0.02fF
C3418 sky130_fd_sc_hd__dfrtn_1_7/a_651_413# DOUT[14] 0.00fF
C3419 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# VDD 0.10fF
C3420 sky130_fd_sc_hd__dfrtn_1_25/a_639_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C3421 sky130_fd_sc_hd__nor3_1_0/a_109_297# VDD 0.00fF
C3422 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_17/a_761_289# 0.01fF
C3423 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_15/A 0.00fF
C3424 sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# sky130_fd_sc_hd__inv_1_32/A 0.01fF
C3425 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# VDD 0.14fF
C3426 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3427 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__mux4_2_0/a_1279_413# 0.00fF
C3428 sky130_fd_sc_hd__dfrtn_1_17/a_805_47# RESET_COUNTERn 0.00fF
C3429 sky130_fd_sc_hd__dfrtn_1_41/a_639_47# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C3430 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__o2111a_2_0/a_386_47# -0.00fF
C3431 sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C3432 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__inv_1_32/A 0.37fF
C3433 RESET_COUNTERn DOUT[14] 0.36fF
C3434 sky130_fd_sc_hd__inv_1_37/A DOUT[10] 0.00fF
C3435 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3436 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C3437 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__mux4_1_0/X 0.06fF
C3438 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C3439 sky130_fd_sc_hd__dfrtn_1_0/a_1270_413# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C3440 sky130_fd_sc_hd__dfrtn_1_19/a_761_289# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C3441 DOUT[4] sky130_fd_sc_hd__dfrtn_1_35/a_1283_21# 0.01fF
C3442 sky130_fd_sc_hd__dfrtn_1_11/a_639_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C3443 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# 0.00fF
C3444 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# 0.00fF
C3445 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# 0.00fF
C3446 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_805_47# 0.00fF
C3447 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_31/a_27_47# 0.03fF
C3448 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C3449 sky130_fd_sc_hd__dfrtn_1_31/a_1270_413# RESET_COUNTERn -0.00fF
C3450 sky130_fd_sc_hd__nor2_1_0/a_109_297# DONE 0.00fF
C3451 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.00fF
C3452 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C3453 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C3454 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_12/a_543_47# 0.00fF
C3455 sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C3456 sky130_fd_sc_hd__dfrtn_1_32/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C3457 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# SEL_CONV_TIME[1] 0.00fF
C3458 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C3459 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_805_47# 0.00fF
C3460 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C3461 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_8/a_761_289# 0.01fF
C3462 CLK_REF sky130_fd_sc_hd__inv_1_28/A 0.18fF
C3463 sky130_fd_sc_hd__dfrtn_1_25/a_651_413# sky130_fd_sc_hd__dfrtn_1_27/a_1217_47# 0.00fF
C3464 sky130_fd_sc_hd__dfrtn_1_20/a_651_413# DOUT[2] 0.00fF
C3465 sky130_fd_sc_hd__inv_1_7/A DOUT[19] 0.01fF
C3466 sky130_fd_sc_hd__inv_1_30/Y DOUT[2] 0.00fF
C3467 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# sky130_fd_sc_hd__dfrtn_1_23/a_543_47# 0.00fF
C3468 sky130_fd_sc_hd__dfrtn_1_22/a_543_47# sky130_fd_sc_hd__dfrtn_1_23/a_193_47# 0.00fF
C3469 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# DOUT[3] 0.02fF
C3470 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_21/a_543_47# 0.00fF
C3471 sky130_fd_sc_hd__dfrtn_1_31/a_448_47# DONE 0.00fF
C3472 sky130_fd_sc_hd__mux4_2_0/a_1279_413# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C3473 sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C3474 sky130_fd_sc_hd__dfrtn_1_38/a_543_47# sky130_fd_sc_hd__inv_1_27/Y 0.00fF
C3475 sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C3476 sky130_fd_sc_hd__inv_1_32/A sky130_fd_sc_hd__inv_1_33/A 0.04fF
C3477 sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C3478 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__inv_1_2/A 0.02fF
C3479 sky130_fd_sc_hd__dfrtn_1_29/a_639_47# SEL_CONV_TIME[0] 0.00fF
C3480 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_33/a_639_47# 0.00fF
C3481 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__dfrtn_1_33/a_1108_47# 0.00fF
C3482 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_33/a_448_47# 0.00fF
C3483 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__dfrtn_1_33/a_651_413# 0.00fF
C3484 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__dfrtn_1_33/a_27_47# 0.00fF
C3485 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__dfrtn_1_33/a_193_47# 0.00fF
C3486 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# 0.00fF
C3487 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__or2_2_0/X 0.01fF
C3488 sky130_fd_sc_hd__dfrtp_1_3/a_761_289# RESET_COUNTERn 0.01fF
C3489 sky130_fd_sc_hd__dfrtn_1_8/a_1462_47# sky130_fd_sc_hd__inv_1_9/Y 0.00fF
C3490 sky130_fd_sc_hd__dfrtn_1_28/a_1217_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C3491 sky130_fd_sc_hd__inv_1_5/A sky130_fd_sc_hd__inv_1_8/A 0.00fF
C3492 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.00fF
C3493 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__o211a_1_1/a_297_297# 0.00fF
C3494 sky130_fd_sc_hd__dfrtn_1_5/a_805_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C3495 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C3496 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# outb 0.00fF
C3497 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3498 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# VDD 0.05fF
C3499 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C3500 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_193_47# 0.00fF
C3501 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_3/a_27_47# 0.00fF
C3502 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C3503 sky130_fd_sc_hd__nor3_1_19/Y SEL_CONV_TIME[3] 0.09fF
C3504 sky130_fd_sc_hd__dfrtn_1_37/a_1462_47# VDD 0.00fF
C3505 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__inv_1_46/Y 0.01fF
C3506 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__inv_1_35/Y 0.00fF
C3507 sky130_fd_sc_hd__dfrtn_1_3/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3508 sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# VDD 0.00fF
C3509 sky130_fd_sc_hd__dfrtn_1_14/a_639_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C3510 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# 0.00fF
C3511 sky130_fd_sc_hd__dfrtp_1_1/a_448_47# sky130_fd_sc_hd__dfrtp_1_2/a_193_47# 0.00fF
C3512 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_2/a_651_413# 0.00fF
C3513 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__dfrtp_1_2/a_27_47# 0.00fF
C3514 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_2/a_448_47# 0.00fF
C3515 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__inv_1_4/A 0.00fF
C3516 sky130_fd_sc_hd__dfrtn_1_34/a_651_413# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C3517 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C3518 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C3519 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__inv_1_53/Y 0.01fF
C3520 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# RESET_COUNTERn 0.00fF
C3521 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C3522 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_805_47# 0.00fF
C3523 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C3524 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C3525 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# 0.00fF
C3526 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_639_47# 0.00fF
C3527 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C3528 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C3529 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C3530 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__inv_1_44/Y 0.54fF
C3531 sky130_fd_sc_hd__dfrtn_1_42/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C3532 sky130_fd_sc_hd__inv_1_44/A sky130_fd_sc_hd__o2111a_2_0/X 0.18fF
C3533 sky130_fd_sc_hd__dfrtn_1_42/a_543_47# VDD 0.05fF
C3534 HEADER_1/a_508_138# sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# 0.00fF
C3535 sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# DOUT[21] 0.00fF
C3536 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# RESET_COUNTERn 0.01fF
C3537 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C3538 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__inv_1_44/A 0.01fF
C3539 sky130_fd_sc_hd__nor3_2_1/a_27_297# DOUT[23] 0.01fF
C3540 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_36/a_543_47# 0.00fF
C3541 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# -0.00fF
C3542 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# -0.00fF
C3543 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# sky130_fd_sc_hd__nor3_1_3/a_109_297# 0.00fF
C3544 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C3545 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C3546 sky130_fd_sc_hd__nor3_1_19/Y SEL_CONV_TIME[2] 0.00fF
C3547 sky130_fd_sc_hd__inv_1_50/Y SEL_CONV_TIME[1] 0.01fF
C3548 sky130_fd_sc_hd__inv_1_38/A sky130_fd_sc_hd__nor3_2_3/C 0.13fF
C3549 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# VDD 0.07fF
C3550 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C3551 sky130_fd_sc_hd__dfrtn_1_9/a_651_413# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C3552 sky130_fd_sc_hd__dfrtn_1_4/a_651_413# VDD 0.01fF
C3553 sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C3554 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# DOUT[11] 0.00fF
C3555 sky130_fd_sc_hd__inv_1_7/Y DOUT[14] 0.00fF
C3556 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.00fF
C3557 sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__dfrtn_1_26/a_761_289# 0.00fF
C3558 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_543_47# 0.00fF
C3559 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__inv_1_31/A 0.00fF
C3560 sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# DOUT[3] 0.01fF
C3561 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# 0.00fF
C3562 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C3563 VDD sky130_fd_sc_hd__inv_1_26/A 0.41fF
C3564 sky130_fd_sc_hd__dfrtn_1_19/a_805_47# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C3565 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# sky130_fd_sc_hd__dfrtn_1_16/a_805_47# -0.00fF
C3566 sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C3567 sky130_fd_sc_hd__dfrtn_1_8/a_27_47# sky130_fd_sc_hd__dfrtn_1_8/a_761_289# -0.00fF
C3568 sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__inv_1_19/A 0.00fF
C3569 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# DOUT[3] 0.00fF
C3570 DOUT[7] DOUT[3] 0.00fF
C3571 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C3572 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.00fF
C3573 sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C3574 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__dfrtn_1_7/a_761_289# 0.00fF
C3575 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__dfrtn_1_7/a_27_47# 0.00fF
C3576 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# sky130_fd_sc_hd__dfrtn_1_7/a_193_47# 0.00fF
C3577 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_543_47# 0.00fF
C3578 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__nor3_1_4/a_109_297# 0.00fF
C3579 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C3580 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_3/a_1108_47# 0.00fF
C3581 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_0/a_448_47# 0.00fF
C3582 sky130_fd_sc_hd__mux4_2_0/a_193_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C3583 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__dfrtn_1_28/a_651_413# -0.00fF
C3584 sky130_fd_sc_hd__dfrtn_1_28/a_193_47# sky130_fd_sc_hd__dfrtn_1_28/a_448_47# -0.00fF
C3585 sky130_fd_sc_hd__nor3_2_2/a_281_297# sky130_fd_sc_hd__dfrtn_1_16/a_1270_413# 0.00fF
C3586 sky130_fd_sc_hd__dfrtp_1_0/a_1108_47# VDD 0.07fF
C3587 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3588 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C3589 DOUT[16] sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C3590 sky130_fd_sc_hd__inv_1_37/A sky130_fd_sc_hd__nor3_2_2/A 0.20fF
C3591 sky130_fd_sc_hd__dfrtn_1_36/a_193_47# sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C3592 sky130_fd_sc_hd__inv_1_2/A DOUT[7] 0.01fF
C3593 sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C3594 sky130_fd_sc_hd__dfrtp_1_1/a_805_47# sky130_fd_sc_hd__o211a_1_1/a_215_47# 0.00fF
C3595 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# DOUT[20] 0.01fF
C3596 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_3/A 0.29fF
C3597 DOUT[19] sky130_fd_sc_hd__inv_1_6/Y 0.04fF
C3598 sky130_fd_sc_hd__dfrtn_1_22/a_1283_21# RESET_COUNTERn 0.02fF
C3599 sky130_fd_sc_hd__dfrtn_1_39/a_448_47# VDD 0.02fF
C3600 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C3601 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C3602 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C3603 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.01fF
C3604 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# 0.00fF
C3605 sky130_fd_sc_hd__nor3_1_11/a_109_297# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C3606 CLK_REF sky130_fd_sc_hd__dfrtn_1_20/a_193_47# 0.01fF
C3607 sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3608 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C3609 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_3/a_27_47# 0.00fF
C3610 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_10/a_761_289# -0.00fF
C3611 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_3/a_639_47# 0.00fF
C3612 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__dfrtn_1_3/a_651_413# 0.00fF
C3613 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# sky130_fd_sc_hd__dfrtn_1_3/a_193_47# 0.00fF
C3614 sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# sky130_fd_sc_hd__dfrtn_1_3/a_27_47# 0.00fF
C3615 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__dfrtn_1_3/a_1270_413# 0.00fF
C3616 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__dfrtn_1_3/a_805_47# 0.00fF
C3617 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C3618 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__inv_1_33/A 0.05fF
C3619 sky130_fd_sc_hd__inv_1_14/A VDD 0.41fF
C3620 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__nor3_2_3/C 0.06fF
C3621 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C3622 sky130_fd_sc_hd__dfrtn_1_18/a_448_47# VDD 0.01fF
C3623 sky130_fd_sc_hd__inv_1_12/A DOUT[3] 0.00fF
C3624 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C3625 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__o221ai_1_0/a_493_297# 0.00fF
C3626 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__inv_1_5/Y 0.02fF
C3627 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_1462_47# 0.00fF
C3628 sky130_fd_sc_hd__dfrtn_1_41/a_1270_413# DOUT[2] 0.00fF
C3629 DOUT[13] DOUT[1] 0.00fF
C3630 sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C3631 VDD en 0.17fF
C3632 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_12/A 0.21fF
C3633 sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C3634 sky130_fd_sc_hd__dfrtn_1_17/a_761_289# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C3635 sky130_fd_sc_hd__dfrtn_1_17/a_543_47# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.01fF
C3636 HEADER_0/a_508_138# DOUT[14] 0.00fF
C3637 sky130_fd_sc_hd__dfrtn_1_42/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3638 sky130_fd_sc_hd__dfrtn_1_16/a_761_289# RESET_COUNTERn 0.01fF
C3639 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# DOUT[14] 0.00fF
C3640 sky130_fd_sc_hd__dfrtn_1_8/a_543_47# DOUT[21] 0.00fF
C3641 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_3/Y 0.04fF
C3642 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_8/Y 0.01fF
C3643 sky130_fd_sc_hd__dfrtn_1_33/a_1108_47# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.01fF
C3644 sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.00fF
C3645 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3646 VDD sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.05fF
C3647 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_20/a_543_47# -0.00fF
C3648 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_20/a_761_289# -0.00fF
C3649 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_651_413# 0.00fF
C3650 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__dfrtn_1_4/a_761_289# 0.00fF
C3651 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C3652 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C3653 sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C3654 SEL_CONV_TIME[0] RESET_COUNTERn 0.24fF
C3655 sky130_fd_sc_hd__dfrtn_1_41/a_805_47# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C3656 sky130_fd_sc_hd__dfrtn_1_41/a_651_413# sky130_fd_sc_hd__dfrtn_1_38/a_543_47# 0.00fF
C3657 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# sky130_fd_sc_hd__dfrtn_1_38/a_651_413# 0.00fF
C3658 sky130_fd_sc_hd__dfrtn_1_41/a_639_47# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C3659 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C3660 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_639_47# 0.00fF
C3661 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_805_47# 0.00fF
C3662 sky130_fd_sc_hd__dfrtn_1_19/a_761_289# VDD 0.05fF
C3663 sky130_fd_sc_hd__dfrtp_1_3/a_1108_47# DOUT[23] 0.00fF
C3664 sky130_fd_sc_hd__nor3_2_2/a_281_297# RESET_COUNTERn 0.00fF
C3665 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__or2b_1_0/a_301_297# 0.00fF
C3666 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_1/a_761_289# 0.00fF
C3667 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_1/a_448_47# 0.00fF
C3668 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_1/a_651_413# 0.00fF
C3669 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_1/a_193_47# 0.00fF
C3670 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C3671 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C3672 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# 0.00fF
C3673 sky130_fd_sc_hd__o221ai_1_0/a_493_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3674 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# 0.00fF
C3675 sky130_fd_sc_hd__o221ai_1_0/a_213_123# VDD 0.01fF
C3676 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__nor3_2_3/B 0.18fF
C3677 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__mux4_2_0/a_1279_413# 0.00fF
C3678 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_18/a_761_289# 0.01fF
C3679 sky130_fd_sc_hd__mux4_2_0/a_872_316# sky130_fd_sc_hd__inv_1_41/Y 0.01fF
C3680 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__inv_1_32/A 0.00fF
C3681 sky130_fd_sc_hd__dfrtn_1_24/a_651_413# SEL_CONV_TIME[1] 0.00fF
C3682 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# sky130_fd_sc_hd__dfrtn_1_7/a_651_413# -0.00fF
C3683 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C3684 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# sky130_fd_sc_hd__o221ai_1_0/a_493_297# 0.00fF
C3685 sky130_fd_sc_hd__dfrtp_1_3/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3686 sky130_fd_sc_hd__nor3_1_0/a_109_297# DOUT[5] 0.00fF
C3687 sky130_fd_sc_hd__dfrtn_1_33/a_639_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C3688 sky130_fd_sc_hd__dfrtn_1_16/a_805_47# DOUT[15] 0.00fF
C3689 sky130_fd_sc_hd__nor3_1_4/a_193_297# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C3690 sky130_fd_sc_hd__nor3_1_5/a_109_297# DOUT[11] 0.00fF
C3691 sky130_fd_sc_hd__nor3_1_1/a_193_297# DOUT[18] 0.00fF
C3692 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C3693 sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# RESET_COUNTERn 0.02fF
C3694 sky130_fd_sc_hd__dfrtn_1_23/a_805_47# DOUT[21] 0.00fF
C3695 sky130_fd_sc_hd__dfrtn_1_22/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3696 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__or3b_2_0/a_27_47# 0.01fF
C3697 sky130_fd_sc_hd__dfrtn_1_26/a_651_413# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C3698 DOUT[10] DOUT[14] 0.00fF
C3699 sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C3700 sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.00fF
C3701 sky130_fd_sc_hd__inv_1_37/A sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C3702 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__dfrtn_1_7/a_1217_47# 0.00fF
C3703 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# sky130_fd_sc_hd__dfrtn_1_7/a_651_413# 0.00fF
C3704 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__dfrtn_1_7/a_639_47# 0.00fF
C3705 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# 0.00fF
C3706 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# sky130_fd_sc_hd__dfrtn_1_7/a_543_47# 0.00fF
C3707 sky130_fd_sc_hd__dfrtn_1_12/a_805_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C3708 sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# DOUT[20] 0.00fF
C3709 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# RESET_COUNTERn -0.01fF
C3710 sky130_fd_sc_hd__dfrtn_1_7/a_543_47# DOUT[7] 0.00fF
C3711 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C3712 DOUT[4] sky130_fd_sc_hd__dfrtn_1_12/a_805_47# 0.00fF
C3713 sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C3714 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C3715 sky130_fd_sc_hd__dfrtn_1_36/a_1462_47# sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C3716 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# sky130_fd_sc_hd__dfrtn_1_0/a_543_47# -0.00fF
C3717 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# DOUT[6] 0.00fF
C3718 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# DOUT[8] 0.00fF
C3719 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# DOUT[7] 0.00fF
C3720 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# RESET_COUNTERn 0.00fF
C3721 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# DOUT[20] 0.00fF
C3722 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# CLK_REF 0.49fF
C3723 DOUT[20] DOUT[7] 0.36fF
C3724 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__inv_1_14/A 0.01fF
C3725 sky130_fd_sc_hd__dfrtn_1_31/a_639_47# sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C3726 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_277_47# -0.00fF
C3727 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_32/a_805_47# 0.00fF
C3728 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C3729 sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C3730 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.00fF
C3731 sky130_fd_sc_hd__dfrtn_1_27/a_543_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C3732 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__inv_1_48/A 0.00fF
C3733 sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C3734 sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3735 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# 0.00fF
C3736 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__o311a_1_0/a_585_47# 0.00fF
C3737 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.00fF
C3738 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C3739 sky130_fd_sc_hd__dfrtn_1_24/a_448_47# VDD 0.01fF
C3740 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C3741 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# VDD 0.08fF
C3742 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__nor3_2_3/C 0.10fF
C3743 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C3744 sky130_fd_sc_hd__dfrtn_1_11/a_639_47# outb 0.00fF
C3745 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3746 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# SEL_CONV_TIME[0] 0.00fF
C3747 sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3748 sky130_fd_sc_hd__nand3b_1_1/Y sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C3749 sky130_fd_sc_hd__inv_1_26/A sky130_fd_sc_hd__o211a_1_0/X 0.00fF
C3750 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__dfrtn_1_3/a_543_47# 0.00fF
C3751 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_31/a_193_47# 0.06fF
C3752 sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# DOUT[14] 0.00fF
C3753 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_52/Y 0.15fF
C3754 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C3755 sky130_fd_sc_hd__nor3_1_19/Y sky130_fd_sc_hd__or3_1_0/X 0.06fF
C3756 sky130_fd_sc_hd__dfrtn_1_17/a_1270_413# sky130_fd_sc_hd__dfrtn_1_19/a_448_47# 0.00fF
C3757 sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# sky130_fd_sc_hd__dfrtn_1_19/a_639_47# 0.00fF
C3758 sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# sky130_fd_sc_hd__dfrtn_1_19/a_805_47# 0.00fF
C3759 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# SEL_CONV_TIME[1] 0.00fF
C3760 sky130_fd_sc_hd__dfrtn_1_26/a_639_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C3761 sky130_fd_sc_hd__dfrtn_1_8/a_639_47# RESET_COUNTERn 0.00fF
C3762 sky130_fd_sc_hd__dfrtp_1_0/a_1108_47# sky130_fd_sc_hd__o211a_1_0/X 0.00fF
C3763 sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3764 sky130_fd_sc_hd__dfrtn_1_30/a_448_47# SEL_CONV_TIME[1] 0.00fF
C3765 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# DOUT[0] 0.00fF
C3766 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__nor3_1_4/a_109_297# 0.00fF
C3767 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# 0.00fF
C3768 sky130_fd_sc_hd__dfrtn_1_20/a_651_413# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C3769 sky130_fd_sc_hd__o211a_1_1/X sky130_fd_sc_hd__or2_2_0/A 0.00fF
C3770 DOUT[15] lc_out 0.00fF
C3771 sky130_fd_sc_hd__inv_1_11/A sky130_fd_sc_hd__inv_1_8/Y 0.01fF
C3772 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_21/a_639_47# 0.00fF
C3773 sky130_fd_sc_hd__dfrtn_1_23/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3774 sky130_fd_sc_hd__dfrtn_1_32/a_1270_413# sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C3775 DOUT[4] sky130_fd_sc_hd__or3b_2_0/a_27_47# 0.00fF
C3776 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_13/a_651_413# 0.00fF
C3777 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# 0.00fF
C3778 sky130_fd_sc_hd__or3b_2_0/a_472_297# sky130_fd_sc_hd__dfrtn_1_30/a_193_47# 0.00fF
C3779 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3780 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__nor3_1_0/A 0.02fF
C3781 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__nand3b_1_1/Y 0.01fF
C3782 sky130_fd_sc_hd__dfrtn_1_24/a_1270_413# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C3783 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C3784 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__inv_1_33/Y 0.02fF
C3785 sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C3786 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# VDD 0.08fF
C3787 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C3788 sky130_fd_sc_hd__inv_1_13/Y sky130_fd_sc_hd__inv_1_13/A 0.01fF
C3789 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__inv_1_51/Y 0.01fF
C3790 SEL_CONV_TIME[0] SEL_CONV_TIME[3] 0.15fF
C3791 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C3792 VDD sky130_fd_sc_hd__or3b_2_0/X 0.05fF
C3793 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__inv_1_47/Y 0.00fF
C3794 sky130_fd_sc_hd__nor3_2_0/a_27_297# RESET_COUNTERn 0.00fF
C3795 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# VDD 0.17fF
C3796 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__dfrtn_1_1/a_448_47# 0.00fF
C3797 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__o2111a_2_0/X -0.04fF
C3798 sky130_fd_sc_hd__o311a_1_0/a_266_297# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C3799 DOUT[4] sky130_fd_sc_hd__nor3_2_3/C 1.57fF
C3800 outb DOUT[12] 0.05fF
C3801 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C3802 sky130_fd_sc_hd__dfrtn_1_7/a_1462_47# RESET_COUNTERn 0.00fF
C3803 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# 0.00fF
C3804 sky130_fd_sc_hd__dfrtn_1_30/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C3805 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# DOUT[3] 0.01fF
C3806 sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# VDD 0.07fF
C3807 sky130_fd_sc_hd__mux4_2_0/a_288_47# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C3808 sky130_fd_sc_hd__dfrtn_1_4/a_651_413# DOUT[3] 0.00fF
C3809 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__a221oi_4_0/a_471_297# 0.01fF
C3810 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3811 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__inv_1_35/A 0.64fF
C3812 sky130_fd_sc_hd__dfrtn_1_16/a_1108_47# DOUT[23] 0.00fF
C3813 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__nor3_1_4/a_109_297# 0.00fF
C3814 DOUT[4] sky130_fd_sc_hd__dfrtn_1_31/a_193_47# 0.00fF
C3815 sky130_fd_sc_hd__dfrtn_1_30/a_543_47# sky130_fd_sc_hd__dfrtn_1_31/a_193_47# 0.00fF
C3816 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__dfrtn_1_31/a_543_47# 0.00fF
C3817 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C3818 sky130_fd_sc_hd__dfrtn_1_14/a_448_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C3819 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# DOUT[14] 0.00fF
C3820 sky130_fd_sc_hd__dfrtn_1_35/a_193_47# sky130_fd_sc_hd__dfrtn_1_35/a_448_47# -0.00fF
C3821 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__dfrtn_1_35/a_651_413# -0.00fF
C3822 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C3823 sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# CLK_REF 0.00fF
C3824 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__inv_1_14/A 0.00fF
C3825 sky130_fd_sc_hd__dfrtn_1_4/a_651_413# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C3826 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__dfrtn_1_17/a_761_289# 0.00fF
C3827 sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C3828 sky130_fd_sc_hd__dfrtn_1_14/a_639_47# DOUT[17] 0.00fF
C3829 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C3830 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__dfrtn_1_17/a_543_47# 0.00fF
C3831 sky130_fd_sc_hd__o211a_1_1/a_510_47# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C3832 sky130_fd_sc_hd__o211a_1_1/a_215_47# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C3833 SEL_CONV_TIME[1] sky130_fd_sc_hd__inv_1_41/Y 0.02fF
C3834 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# SEL_CONV_TIME[1] 0.00fF
C3835 SEL_CONV_TIME[0] SEL_CONV_TIME[2] 0.03fF
C3836 DOUT[15] sky130_fd_sc_hd__nor3_2_3/B 0.52fF
C3837 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C3838 sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__o211a_1_0/a_79_21# 0.06fF
C3839 sky130_fd_sc_hd__dfrtn_1_16/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3840 sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# VDD -0.00fF
C3841 sky130_fd_sc_hd__dfrtn_1_8/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3842 sky130_fd_sc_hd__dfrtn_1_5/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3843 sky130_fd_sc_hd__o211a_1_0/a_79_21# sky130_fd_sc_hd__o211a_1_0/a_215_47# -0.00fF
C3844 sky130_fd_sc_hd__dfrtn_1_36/a_651_413# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C3845 sky130_fd_sc_hd__or3_1_0/a_111_297# sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C3846 sky130_fd_sc_hd__nor3_1_1/a_193_297# DOUT[22] 0.00fF
C3847 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C3848 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__nor3_1_3/a_193_297# 0.00fF
C3849 sky130_fd_sc_hd__nor3_1_19/Y sky130_fd_sc_hd__inv_1_53/A 0.00fF
C3850 sky130_fd_sc_hd__inv_1_19/A sky130_fd_sc_hd__inv_1_22/A 0.00fF
C3851 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# 0.00fF
C3852 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__dfrtn_1_11/a_193_47# 0.00fF
C3853 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_11/a_543_47# 0.00fF
C3854 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# sky130_fd_sc_hd__dfrtn_1_11/a_761_289# 0.00fF
C3855 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C3856 sky130_fd_sc_hd__o211a_1_1/a_215_47# VDD 0.00fF
C3857 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3858 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C3859 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C3860 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_12/a_1270_413# 0.00fF
C3861 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C3862 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# 0.00fF
C3863 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# 0.00fF
C3864 DOUT[4] sky130_fd_sc_hd__dfrtn_1_32/a_448_47# 0.01fF
C3865 sky130_fd_sc_hd__o2111a_2_0/a_386_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C3866 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_1/a_193_47# -0.32fF
C3867 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C3868 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# sky130_fd_sc_hd__inv_1_6/A 0.25fF
C3869 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C3870 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# 0.00fF
C3871 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C3872 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# 0.00fF
C3873 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# 0.01fF
C3874 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_17/a_651_413# 0.00fF
C3875 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__dfrtn_1_17/a_761_289# 0.00fF
C3876 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_639_47# 0.00fF
C3877 sky130_fd_sc_hd__dfrtp_1_2/a_639_47# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C3878 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__dfrtn_1_17/a_448_47# 0.00fF
C3879 sky130_fd_sc_hd__nor3_2_2/A DOUT[14] 0.00fF
C3880 sky130_fd_sc_hd__dfrtn_1_12/a_639_47# sky130_fd_sc_hd__dfrtn_1_14/a_27_47# 0.00fF
C3881 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_14/a_639_47# 0.00fF
C3882 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# 0.00fF
C3883 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__dfrtn_1_14/a_543_47# 0.00fF
C3884 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C3885 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_14/a_543_47# 0.00fF
C3886 sky130_fd_sc_hd__dfrtn_1_28/a_193_47# sky130_fd_sc_hd__or3_1_0/C 0.01fF
C3887 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__dfrtn_1_42/a_448_47# 0.00fF
C3888 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# VDD 0.17fF
C3889 sky130_fd_sc_hd__o211a_1_0/a_79_21# sky130_fd_sc_hd__or2_2_0/B 0.01fF
C3890 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C3891 VDD VIN 2.76fF
C3892 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C3893 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# DOUT[14] 0.00fF
C3894 sky130_fd_sc_hd__nor3_1_12/a_109_297# outb 0.00fF
C3895 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# VDD 0.12fF
C3896 sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C3897 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# VDD 0.00fF
C3898 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__dfrtn_1_30/a_193_47# 0.00fF
C3899 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__dfrtn_1_30/a_27_47# 0.00fF
C3900 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# sky130_fd_sc_hd__o221ai_1_0/a_493_297# 0.00fF
C3901 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C3902 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__inv_1_40/Y 0.14fF
C3903 sky130_fd_sc_hd__dfrtn_1_28/a_193_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C3904 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C3905 sky130_fd_sc_hd__dfrtn_1_7/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3906 sky130_fd_sc_hd__dfrtn_1_16/a_1283_21# sky130_fd_sc_hd__inv_1_26/A 0.00fF
C3907 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3908 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# VDD 0.00fF
C3909 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# DOUT[21] 0.00fF
C3910 sky130_fd_sc_hd__nor3_2_1/a_27_297# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C3911 sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# sky130_fd_sc_hd__dfrtn_1_23/a_448_47# 0.00fF
C3912 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C3913 sky130_fd_sc_hd__dfrtn_1_37/a_1270_413# RESET_COUNTERn 0.00fF
C3914 sky130_fd_sc_hd__dfrtn_1_32/a_543_47# sky130_fd_sc_hd__inv_1_36/A 0.01fF
C3915 sky130_fd_sc_hd__nor3_1_1/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3916 SEL_CONV_TIME[1] sky130_fd_sc_hd__inv_1_49/A 0.04fF
C3917 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C3918 DOUT[9] sky130_fd_sc_hd__dfrtn_1_6/a_193_47# 0.00fF
C3919 sky130_fd_sc_hd__dfrtn_1_33/a_1217_47# VDD 0.00fF
C3920 sky130_fd_sc_hd__dfrtn_1_33/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3921 sky130_fd_sc_hd__dfrtn_1_3/a_651_413# RESET_COUNTERn 0.00fF
C3922 sky130_fd_sc_hd__dfrtn_1_31/a_805_47# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C3923 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__inv_1_43/A 0.02fF
C3924 outb sky130_fd_sc_hd__nor3_2_3/C 1.57fF
C3925 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C3926 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# HEADER_0/a_508_138# 0.00fF
C3927 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C3928 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# VDD 0.10fF
C3929 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3930 sky130_fd_sc_hd__dfrtn_1_20/a_1217_47# sky130_fd_sc_hd__inv_1_35/A 0.00fF
C3931 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C3932 sky130_fd_sc_hd__dfrtn_1_34/a_543_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C3933 sky130_fd_sc_hd__dfrtn_1_0/a_543_47# sky130_fd_sc_hd__inv_1_15/A 0.01fF
C3934 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C3935 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C3936 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# HEADER_0/a_508_138# 0.00fF
C3937 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__or2_2_0/B 0.03fF
C3938 DOUT[13] sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# 0.00fF
C3939 sky130_fd_sc_hd__dfrtn_1_0/a_448_47# DOUT[17] 0.00fF
C3940 sky130_fd_sc_hd__dfrtn_1_17/a_543_47# sky130_fd_sc_hd__inv_1_28/A 0.01fF
C3941 sky130_fd_sc_hd__nor3_1_3/a_109_297# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C3942 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# DOUT[6] 0.00fF
C3943 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# DOUT[8] 0.00fF
C3944 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# RESET_COUNTERn 0.16fF
C3945 sky130_fd_sc_hd__dfrtn_1_24/a_805_47# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C3946 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# sky130_fd_sc_hd__dfrtn_1_29/a_761_289# 0.00fF
C3947 sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C3948 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# sky130_fd_sc_hd__dfrtn_1_29/a_639_47# 0.00fF
C3949 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_29/a_805_47# 0.00fF
C3950 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# 0.00fF
C3951 DOUT[11] sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C3952 sky130_fd_sc_hd__dfrtn_1_4/a_543_47# RESET_COUNTERn 0.01fF
C3953 sky130_fd_sc_hd__nor3_2_0/A sky130_fd_sc_hd__inv_1_8/Y 0.02fF
C3954 sky130_fd_sc_hd__dfrtn_1_38/a_639_47# VDD 0.00fF
C3955 sky130_fd_sc_hd__dfrtn_1_33/a_651_413# sky130_fd_sc_hd__inv_1_45/A 0.00fF
C3956 sky130_fd_sc_hd__nor3_1_5/a_193_297# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C3957 sky130_fd_sc_hd__dfrtn_1_21/a_805_47# RESET_COUNTERn 0.00fF
C3958 sky130_fd_sc_hd__nor3_1_20/a_109_297# DOUT[1] 0.00fF
C3959 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__dfrtn_1_11/a_1462_47# 0.00fF
C3960 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# sky130_fd_sc_hd__dfrtn_1_11/a_1270_413# 0.00fF
C3961 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__dfrtn_1_11/a_639_47# 0.00fF
C3962 sky130_fd_sc_hd__dfrtn_1_10/a_1217_47# sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# 0.00fF
C3963 sky130_fd_sc_hd__dfrtn_1_10/a_805_47# sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# 0.00fF
C3964 sky130_fd_sc_hd__inv_1_28/A sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3965 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C3966 sky130_fd_sc_hd__inv_1_4/Y DOUT[14] 0.35fF
C3967 sky130_fd_sc_hd__dfrtn_1_42/a_651_413# DOUT[15] 0.00fF
C3968 sky130_fd_sc_hd__inv_1_0/A VDD 0.58fF
C3969 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C3970 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# -0.00fF
C3971 sky130_fd_sc_hd__dfrtn_1_7/a_1217_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C3972 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_40/a_27_47# 0.00fF
C3973 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# VDD 0.08fF
C3974 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# 0.00fF
C3975 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# -0.00fF
C3976 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__dfrtn_1_0/a_761_289# 0.00fF
C3977 sky130_fd_sc_hd__dfrtn_1_12/a_761_289# sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# 0.00fF
C3978 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# 0.00fF
C3979 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# sky130_fd_sc_hd__dfrtn_1_0/a_193_47# 0.00fF
C3980 sky130_fd_sc_hd__or2_2_0/a_121_297# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C3981 sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# VDD 0.00fF
C3982 sky130_fd_sc_hd__dfrtn_1_26/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3983 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_0/a_27_47# 0.00fF
C3984 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# DOUT[3] 0.00fF
C3985 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# RESET_COUNTERn 0.02fF
C3986 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__inv_1_45/Y 0.01fF
C3987 sky130_fd_sc_hd__dfrtn_1_34/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C3988 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C3989 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# -0.00fF
C3990 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# -0.00fF
C3991 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# sky130_fd_sc_hd__dfrtn_1_41/a_543_47# -0.00fF
C3992 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C3993 sky130_fd_sc_hd__dfrtn_1_34/a_1462_47# VDD 0.00fF
C3994 sky130_fd_sc_hd__nor3_1_11/a_193_297# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C3995 sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C3996 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# 0.00fF
C3997 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# 0.00fF
C3998 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_8/a_448_47# 0.00fF
C3999 SLC_0/a_1235_416# DOUT[15] 0.00fF
C4000 sky130_fd_sc_hd__dfrtn_1_23/a_1217_47# sky130_fd_sc_hd__inv_1_40/Y 0.00fF
C4001 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C4002 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_639_47# -0.00fF
C4003 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__inv_1_2/A 0.02fF
C4004 sky130_fd_sc_hd__dfrtn_1_21/a_448_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C4005 sky130_fd_sc_hd__dfrtn_1_39/a_761_289# RESET_COUNTERn 0.00fF
C4006 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__inv_1_39/Y 0.55fF
C4007 DOUT[13] sky130_fd_sc_hd__dfrtn_1_32/a_193_47# 0.00fF
C4008 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_21/a_1270_413# 0.00fF
C4009 sky130_fd_sc_hd__dfrtn_1_25/a_639_47# RESET_COUNTERn 0.00fF
C4010 VDD sky130_fd_sc_hd__inv_1_1/A 0.46fF
C4011 sky130_fd_sc_hd__dfrtp_1_3/a_1108_47# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C4012 sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C4013 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# sky130_fd_sc_hd__inv_1_32/Y 0.00fF
C4014 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C4015 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C4016 sky130_fd_sc_hd__dfrtp_1_3/a_448_47# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.00fF
C4017 sky130_fd_sc_hd__nor3_1_15/a_193_297# DOUT[4] 0.00fF
C4018 sky130_fd_sc_hd__dfrtn_1_18/a_761_289# RESET_COUNTERn 0.00fF
C4019 sky130_fd_sc_hd__dfrtp_1_0/a_639_47# DOUT[15] 0.00fF
C4020 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_26/a_651_413# 0.00fF
C4021 DOUT[15] DOUT[0] 0.00fF
C4022 sky130_fd_sc_hd__inv_1_40/Y RESET_COUNTERn 0.05fF
C4023 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C4024 sky130_fd_sc_hd__or3_1_0/a_111_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4025 en DOUT[20] 0.02fF
C4026 sky130_fd_sc_hd__dfrtn_1_7/a_1462_47# HEADER_0/a_508_138# 0.00fF
C4027 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C4028 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C4029 sky130_fd_sc_hd__or3_1_0/X SEL_CONV_TIME[0] 0.02fF
C4030 sky130_fd_sc_hd__dfrtn_1_28/a_448_47# SEL_CONV_TIME[1] 0.00fF
C4031 sky130_fd_sc_hd__dfrtn_1_42/a_805_47# RESET_COUNTERn 0.00fF
C4032 sky130_fd_sc_hd__mux4_2_0/a_397_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C4033 sky130_fd_sc_hd__dfrtn_1_37/a_1270_413# SEL_CONV_TIME[3] 0.00fF
C4034 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# DOUT[3] 0.15fF
C4035 sky130_fd_sc_hd__dfrtn_1_11/a_1270_413# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C4036 sky130_fd_sc_hd__mux4_2_0/a_872_316# sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.00fF
C4037 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__o311a_1_0/a_266_47# 0.00fF
C4038 sky130_fd_sc_hd__inv_1_3/Y DOUT[7] 0.01fF
C4039 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_10/a_805_47# 0.00fF
C4040 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C4041 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtp_1_3/a_651_413# 0.00fF
C4042 sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C4043 sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C4044 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C4045 CLK_REF sky130_fd_sc_hd__dfrtn_1_17/a_761_289# 0.01fF
C4046 sky130_fd_sc_hd__dfrtn_1_22/a_1283_21# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C4047 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__inv_1_2/A 0.02fF
C4048 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# RESET_COUNTERn 0.00fF
C4049 sky130_fd_sc_hd__dfrtn_1_24/a_1270_413# SEL_CONV_TIME[0] 0.00fF
C4050 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__nor3_2_3/A 0.13fF
C4051 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__inv_1_12/A 0.01fF
C4052 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4053 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__o2111a_2_0/a_80_21# 0.01fF
C4054 sky130_fd_sc_hd__or2b_1_0/a_301_297# sky130_fd_sc_hd__dfrtn_1_34/a_448_47# 0.00fF
C4055 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__nor3_1_3/a_109_297# 0.00fF
C4056 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# -0.03fF
C4057 sky130_fd_sc_hd__dfrtn_1_31/a_639_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C4058 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_761_289# 0.00fF
C4059 sky130_fd_sc_hd__dfrtn_1_35/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C4060 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_25/a_761_289# -0.00fF
C4061 DOUT[13] sky130_fd_sc_hd__dfrtn_1_31/a_651_413# 0.00fF
C4062 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# 0.00fF
C4063 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# 0.01fF
C4064 sky130_fd_sc_hd__inv_1_27/A DOUT[2] 0.27fF
C4065 sky130_fd_sc_hd__dfrtn_1_37/a_1270_413# SEL_CONV_TIME[2] 0.00fF
C4066 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_29/a_651_413# 0.00fF
C4067 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_7/Y 0.01fF
C4068 sky130_fd_sc_hd__dfrtn_1_28/a_1108_47# VDD 0.07fF
C4069 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C4070 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# sky130_fd_sc_hd__inv_1_39/Y 0.00fF
C4071 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# -0.00fF
C4072 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_448_47# -0.00fF
C4073 sky130_fd_sc_hd__dfrtn_1_4/a_543_47# sky130_fd_sc_hd__inv_1_7/Y 0.01fF
C4074 sky130_fd_sc_hd__dfrtn_1_14/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4075 sky130_fd_sc_hd__dfrtn_1_25/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C4076 sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# VDD 0.00fF
C4077 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_12/A 0.00fF
C4078 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_37/a_27_47# 0.05fF
C4079 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# sky130_fd_sc_hd__inv_1_12/A 0.68fF
C4080 sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C4081 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_21/a_761_289# 0.01fF
C4082 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C4083 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__nor3_2_3/B 0.25fF
C4084 sky130_fd_sc_hd__dfrtn_1_16/a_761_289# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C4085 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_0/a_1217_47# 0.00fF
C4086 sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# DOUT[3] 0.00fF
C4087 sky130_fd_sc_hd__nor3_1_10/a_193_297# sky130_fd_sc_hd__inv_1_4/A 0.00fF
C4088 sky130_fd_sc_hd__dfrtp_1_0/a_1462_47# RESET_COUNTERn 0.00fF
C4089 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__dfrtn_1_29/a_448_47# 0.00fF
C4090 DOUT[9] sky130_fd_sc_hd__nor3_1_0/a_193_297# 0.00fF
C4091 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C4092 sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C4093 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__inv_1_37/A 0.01fF
C4094 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C4095 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_38/a_761_289# 0.01fF
C4096 DOUT[9] sky130_fd_sc_hd__dfrtn_1_3/a_193_47# 0.00fF
C4097 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C4098 sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C4099 sky130_fd_sc_hd__nor3_2_2/a_281_297# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C4100 sky130_fd_sc_hd__dfrtn_1_24/a_805_47# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C4101 sky130_fd_sc_hd__inv_1_36/Y RESET_COUNTERn 0.00fF
C4102 sky130_fd_sc_hd__dfrtn_1_22/a_1217_47# sky130_fd_sc_hd__inv_1_39/Y 0.00fF
C4103 sky130_fd_sc_hd__dfrtn_1_20/a_543_47# VDD 0.04fF
C4104 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C4105 sky130_fd_sc_hd__dfrtn_1_42/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4106 sky130_fd_sc_hd__dfrtn_1_24/a_651_413# DOUT[21] 0.01fF
C4107 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# RESET_COUNTERn 0.00fF
C4108 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# DOUT[20] 0.00fF
C4109 sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# sky130_fd_sc_hd__inv_1_42/A 0.01fF
C4110 VDD sky130_fd_sc_hd__inv_1_11/A 0.34fF
C4111 CLK_REF sky130_fd_sc_hd__nor3_2_1/a_27_297# 0.00fF
C4112 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__o2111a_2_0/a_566_47# 0.00fF
C4113 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__o2111a_2_0/a_458_47# 0.00fF
C4114 sky130_fd_sc_hd__inv_1_30/A RESET_COUNTERn 0.12fF
C4115 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__dfrtn_1_25/a_651_413# 0.00fF
C4116 DOUT[1] sky130_fd_sc_hd__dfrtn_1_36/a_543_47# 0.00fF
C4117 sky130_fd_sc_hd__inv_1_53/A SEL_CONV_TIME[0] 0.01fF
C4118 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_13/Y 0.07fF
C4119 VIN DOUT[3] 0.16fF
C4120 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.09fF
C4121 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4122 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# DOUT[2] 0.01fF
C4123 sky130_fd_sc_hd__dfrtn_1_22/a_1108_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C4124 sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4125 sky130_fd_sc_hd__dfrtn_1_42/a_193_47# sky130_fd_sc_hd__dfrtn_1_42/a_543_47# -0.00fF
C4126 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# -0.00fF
C4127 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__inv_1_50/A 0.00fF
C4128 sky130_fd_sc_hd__dfrtn_1_30/a_651_413# SEL_CONV_TIME[0] 0.01fF
C4129 sky130_fd_sc_hd__dfrtn_1_25/a_639_47# SEL_CONV_TIME[3] 0.00fF
C4130 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__dfrtn_1_7/a_448_47# 0.00fF
C4131 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__nor3_2_3/B 0.03fF
C4132 sky130_fd_sc_hd__nor3_1_14/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4133 sky130_fd_sc_hd__inv_1_2/A VIN 0.13fF
C4134 sky130_fd_sc_hd__inv_1_34/Y sky130_fd_sc_hd__inv_1_28/Y 0.01fF
C4135 sky130_fd_sc_hd__mux4_1_0/a_923_363# VDD 0.00fF
C4136 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4137 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# DOUT[3] 0.00fF
C4138 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C4139 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__inv_1_33/A 0.01fF
C4140 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4141 sky130_fd_sc_hd__dfrtn_1_10/a_1270_413# VDD 0.00fF
C4142 sky130_fd_sc_hd__dfrtn_1_9/a_805_47# RESET_COUNTERn 0.00fF
C4143 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C4144 sky130_fd_sc_hd__dfrtn_1_11/a_761_289# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C4145 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# 0.00fF
C4146 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# sky130_fd_sc_hd__dfrtn_1_15/a_27_47# 0.00fF
C4147 sky130_fd_sc_hd__dfrtp_1_0/a_1283_21# DOUT[23] 0.00fF
C4148 sky130_fd_sc_hd__dfrtn_1_24/a_651_413# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C4149 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C4150 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C4151 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_761_289# -0.00fF
C4152 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__nor3_1_19/Y 0.01fF
C4153 sky130_fd_sc_hd__dfrtn_1_19/a_639_47# RESET_COUNTERn 0.00fF
C4154 sky130_fd_sc_hd__nor3_1_8/a_109_297# DOUT[8] 0.00fF
C4155 sky130_fd_sc_hd__nor3_1_8/a_193_297# DOUT[7] 0.00fF
C4156 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C4157 sky130_fd_sc_hd__nor3_1_4/a_193_297# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C4158 sky130_fd_sc_hd__mux4_2_0/a_397_47# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C4159 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_11/a_193_47# 0.00fF
C4160 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C4161 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# sky130_fd_sc_hd__inv_1_49/A 0.02fF
C4162 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# SEL_CONV_TIME[0] 0.00fF
C4163 sky130_fd_sc_hd__mux4_2_0/a_600_345# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C4164 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_448_47# -0.00fF
C4165 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# -0.00fF
C4166 sky130_fd_sc_hd__inv_1_39/A sky130_fd_sc_hd__inv_1_40/A 0.01fF
C4167 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# DOUT[6] 0.00fF
C4168 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# DOUT[20] 0.00fF
C4169 sky130_fd_sc_hd__dfrtp_1_0/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4170 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_4/a_651_413# 0.00fF
C4171 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__dfrtn_1_4/a_448_47# 0.00fF
C4172 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C4173 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C4174 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C4175 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C4176 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C4177 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C4178 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C4179 sky130_fd_sc_hd__dfrtn_1_39/a_761_289# SEL_CONV_TIME[2] 0.01fF
C4180 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C4181 sky130_fd_sc_hd__dfrtn_1_35/a_1462_47# DOUT[16] 0.00fF
C4182 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_40/a_1270_413# 0.00fF
C4183 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__inv_1_45/A 0.00fF
C4184 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C4185 sky130_fd_sc_hd__dfrtn_1_27/a_448_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C4186 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C4187 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C4188 sky130_fd_sc_hd__dfrtn_1_12/a_1270_413# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C4189 sky130_fd_sc_hd__dfrtn_1_0/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4190 sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C4191 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# 0.00fF
C4192 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C4193 sky130_fd_sc_hd__dfrtn_1_35/a_1108_47# VDD 0.07fF
C4194 sky130_fd_sc_hd__dfrtn_1_0/a_639_47# VDD 0.00fF
C4195 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# sky130_fd_sc_hd__inv_1_15/A 0.02fF
C4196 sky130_fd_sc_hd__o311a_1_0/a_81_21# SEL_CONV_TIME[1] 0.01fF
C4197 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# RESET_COUNTERn 0.31fF
C4198 sky130_fd_sc_hd__inv_1_42/Y SEL_CONV_TIME[0] 0.35fF
C4199 sky130_fd_sc_hd__dfrtn_1_26/a_761_289# SEL_CONV_TIME[0] 0.00fF
C4200 sky130_fd_sc_hd__dfrtn_1_12/a_1270_413# DOUT[17] 0.00fF
C4201 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C4202 sky130_fd_sc_hd__dfrtn_1_3/a_639_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C4203 sky130_fd_sc_hd__mux4_2_0/a_193_369# SEL_CONV_TIME[1] -0.00fF
C4204 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# DOUT[19] 0.00fF
C4205 sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# sky130_fd_sc_hd__or3_1_0/C 0.02fF
C4206 sky130_fd_sc_hd__dfrtn_1_34/a_543_47# SEL_CONV_TIME[0] 0.01fF
C4207 sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C4208 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# VDD 0.05fF
C4209 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.03fF
C4210 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# 0.00fF
C4211 sky130_fd_sc_hd__inv_1_42/A sky130_fd_sc_hd__inv_1_48/A 0.00fF
C4212 sky130_fd_sc_hd__inv_1_50/A DOUT[4] 0.43fF
C4213 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C4214 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C4215 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_30/a_543_47# 0.00fF
C4216 sky130_fd_sc_hd__dfrtn_1_39/a_805_47# sky130_fd_sc_hd__inv_1_32/Y 0.00fF
C4217 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C4218 sky130_fd_sc_hd__or3_1_0/a_183_297# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C4219 sky130_fd_sc_hd__inv_1_54/Y DOUT[2] 0.04fF
C4220 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_448_47# -0.00fF
C4221 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# -0.00fF
C4222 sky130_fd_sc_hd__dfrtn_1_21/a_448_47# VDD 0.01fF
C4223 sky130_fd_sc_hd__dfrtp_1_0/a_761_289# SLC_0/a_438_293# 0.00fF
C4224 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# SLC_0/a_919_243# 0.00fF
C4225 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# SLC_0/a_264_22# 0.01fF
C4226 sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# RESET_COUNTERn 0.00fF
C4227 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# sky130_fd_sc_hd__inv_1_26/A 0.00fF
C4228 sky130_fd_sc_hd__inv_1_45/Y SEL_CONV_TIME[1] 0.00fF
C4229 sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4230 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__nand3b_1_0/a_53_93# 0.00fF
C4231 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# SEL_CONV_TIME[1] 0.00fF
C4232 sky130_fd_sc_hd__dfrtn_1_42/a_1108_47# sky130_fd_sc_hd__inv_1_40/Y 0.00fF
C4233 VDD sky130_fd_sc_hd__inv_1_39/A 0.38fF
C4234 CLK_REF sky130_fd_sc_hd__dfrtp_1_3/a_1108_47# 0.01fF
C4235 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__dfrtn_1_24/a_27_47# 0.00fF
C4236 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# 0.00fF
C4237 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# 0.00fF
C4238 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C4239 sky130_fd_sc_hd__dfrtn_1_8/a_761_289# outb 0.00fF
C4240 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_44/A 0.21fF
C4241 DOUT[15] DOUT[2] 0.08fF
C4242 sky130_fd_sc_hd__inv_1_0/A DOUT[5] 0.00fF
C4243 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_12/a_651_413# -0.00fF
C4244 sky130_fd_sc_hd__nand3b_1_0/a_316_47# SEL_CONV_TIME[1] 0.00fF
C4245 sky130_fd_sc_hd__dfrtn_1_16/a_1217_47# DOUT[2] 0.00fF
C4246 sky130_fd_sc_hd__inv_1_36/A DOUT[21] 0.02fF
C4247 DOUT[9] sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# 0.00fF
C4248 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# 0.00fF
C4249 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__dfrtn_1_13/a_543_47# 0.00fF
C4250 sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# 0.00fF
C4251 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# sky130_fd_sc_hd__dfrtn_1_13/a_761_289# 0.00fF
C4252 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_12/a_761_289# 0.00fF
C4253 sky130_fd_sc_hd__dfrtn_1_7/a_543_47# VIN 0.04fF
C4254 DOUT[9] sky130_fd_sc_hd__dfrtn_1_4/a_1270_413# 0.00fF
C4255 sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# DOUT[11] 0.00fF
C4256 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__inv_1_5/Y 0.01fF
C4257 sky130_fd_sc_hd__o211a_1_1/X RESET_COUNTERn 0.00fF
C4258 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__dfrtp_1_0/a_651_413# -0.00fF
C4259 sky130_fd_sc_hd__mux4_2_0/a_27_47# VDD 0.12fF
C4260 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# out 0.01fF
C4261 sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C4262 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# VIN 0.00fF
C4263 sky130_fd_sc_hd__inv_1_1/A DOUT[3] 0.14fF
C4264 sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C4265 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__nor3_2_1/a_281_297# 0.00fF
C4266 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__nor3_2_1/a_27_297# 0.00fF
C4267 VIN DOUT[20] 0.11fF
C4268 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C4269 sky130_fd_sc_hd__inv_1_6/A sky130_fd_sc_hd__inv_1_2/Y 0.01fF
C4270 sky130_fd_sc_hd__nor3_1_13/a_193_297# RESET_COUNTERn 0.00fF
C4271 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__inv_1_38/Y 0.06fF
C4272 sky130_fd_sc_hd__inv_1_41/Y DOUT[21] 0.00fF
C4273 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# DOUT[21] 0.00fF
C4274 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__inv_1_23/A 0.01fF
C4275 sky130_fd_sc_hd__dfrtn_1_5/a_805_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C4276 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# RESET_COUNTERn 0.03fF
C4277 sky130_fd_sc_hd__nor3_1_0/a_109_297# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C4278 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_11/a_1462_47# 0.00fF
C4279 VDD sky130_fd_sc_hd__inv_1_35/A 0.54fF
C4280 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_1/A 0.00fF
C4281 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# VDD 0.09fF
C4282 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# DOUT[6] 0.00fF
C4283 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# RESET_COUNTERn 0.00fF
C4284 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C4285 sky130_fd_sc_hd__dfrtn_1_39/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_639_47# -0.00fF
C4286 sky130_fd_sc_hd__inv_1_1/A DOUT[5] 0.01fF
C4287 sky130_fd_sc_hd__inv_1_19/A DOUT[12] 0.00fF
C4288 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C4289 sky130_fd_sc_hd__nand3b_1_0/a_232_47# VDD 0.00fF
C4290 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# 0.00fF
C4291 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C4292 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__inv_1_45/A 0.00fF
C4293 sky130_fd_sc_hd__o311a_1_0/a_266_297# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C4294 sky130_fd_sc_hd__dfrtn_1_39/a_448_47# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C4295 sky130_fd_sc_hd__dfrtn_1_33/a_651_413# RESET_COUNTERn 0.00fF
C4296 DOUT[1] sky130_fd_sc_hd__dfrtn_1_32/a_805_47# 0.00fF
C4297 sky130_fd_sc_hd__dfrtn_1_7/a_651_413# DOUT[19] 0.00fF
C4298 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# 0.01fF
C4299 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__mux4_2_0/a_1279_413# 0.00fF
C4300 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__mux4_2_0/a_1064_47# 0.00fF
C4301 VDD sky130_fd_sc_hd__nor3_2_0/A 0.57fF
C4302 sky130_fd_sc_hd__mux4_2_0/a_288_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C4303 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4304 sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# RESET_COUNTERn 0.00fF
C4305 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# 0.01fF
C4306 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C4307 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_805_47# 0.00fF
C4308 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C4309 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.00fF
C4310 sky130_fd_sc_hd__inv_1_41/Y sky130_fd_sc_hd__o311a_1_0/A3 0.09fF
C4311 SEL_CONV_TIME[1] sky130_fd_sc_hd__or3_1_0/C 0.11fF
C4312 sky130_fd_sc_hd__mux4_2_0/a_1281_47# SEL_CONV_TIME[1] 0.00fF
C4313 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# RESET_COUNTERn 0.05fF
C4314 VDD DOUT[17] 2.07fF
C4315 DOUT[19] RESET_COUNTERn 0.05fF
C4316 sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C4317 sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4318 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C4319 sky130_fd_sc_hd__nor3_1_16/a_193_297# sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C4320 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__inv_1_11/A 0.01fF
C4321 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C4322 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# sky130_fd_sc_hd__inv_1_47/A 0.01fF
C4323 sky130_fd_sc_hd__or2b_1_0/X SEL_CONV_TIME[1] 0.08fF
C4324 DOUT[1] sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C4325 sky130_fd_sc_hd__dfrtn_1_30/a_805_47# DONE 0.00fF
C4326 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__or2_2_0/X 0.00fF
C4327 sky130_fd_sc_hd__dfrtp_1_0/a_1217_47# SLC_0/a_919_243# 0.00fF
C4328 sky130_fd_sc_hd__dfrtp_1_0/a_1462_47# SLC_0/a_264_22# 0.00fF
C4329 sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# RESET_COUNTERn 0.03fF
C4330 sky130_fd_sc_hd__dfrtn_1_14/a_651_413# DOUT[18] 0.00fF
C4331 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__o211a_1_1/a_297_297# 0.00fF
C4332 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C4333 sky130_fd_sc_hd__inv_1_49/A DOUT[21] 0.00fF
C4334 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C4335 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C4336 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.00fF
C4337 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C4338 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C4339 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# 0.00fF
C4340 sky130_fd_sc_hd__nor3_2_3/a_281_297# RESET_COUNTERn 0.02fF
C4341 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# VDD 0.15fF
C4342 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C4343 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_10/a_1270_413# 0.00fF
C4344 sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C4345 sky130_fd_sc_hd__dfrtn_1_17/a_193_47# sky130_fd_sc_hd__inv_1_28/Y 0.07fF
C4346 outb sky130_fd_sc_hd__inv_1_12/A 0.00fF
C4347 sky130_fd_sc_hd__mux4_2_0/a_1279_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4348 sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C4349 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C4350 sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# DOUT[5] 0.00fF
C4351 sky130_fd_sc_hd__mux4_2_0/a_1064_47# VDD 0.00fF
C4352 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__inv_1_33/A 0.20fF
C4353 sky130_fd_sc_hd__dfrtn_1_9/a_543_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C4354 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# -0.00fF
C4355 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# -0.00fF
C4356 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# DOUT[14] 0.00fF
C4357 sky130_fd_sc_hd__nor3_1_6/a_109_297# DOUT[11] 0.00fF
C4358 sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# sky130_fd_sc_hd__inv_1_33/A 0.03fF
C4359 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__o311a_1_0/a_368_297# 0.00fF
C4360 sky130_fd_sc_hd__dfrtn_1_26/a_651_413# RESET_COUNTERn 0.00fF
C4361 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_2/a_651_413# 0.00fF
C4362 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_34/a_27_47# 0.00fF
C4363 sky130_fd_sc_hd__dfrtn_1_37/a_1270_413# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C4364 VDD sky130_fd_sc_hd__inv_1_28/Y 0.48fF
C4365 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# sky130_fd_sc_hd__dfrtp_1_3/a_761_289# 0.00fF
C4366 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C4367 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__dfrtp_1_3/a_543_47# 0.00fF
C4368 sky130_fd_sc_hd__dfrtp_1_1/a_448_47# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C4369 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_3/a_448_47# 0.00fF
C4370 sky130_fd_sc_hd__dfrtn_1_16/a_448_47# sky130_fd_sc_hd__nor3_2_3/A 0.01fF
C4371 sky130_fd_sc_hd__dfrtn_1_11/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4372 sky130_fd_sc_hd__dfrtn_1_34/a_1270_413# RESET_COUNTERn 0.00fF
C4373 sky130_fd_sc_hd__dfrtn_1_33/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4374 sky130_fd_sc_hd__dfrtn_1_11/a_805_47# VDD 0.00fF
C4375 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_21/a_1217_47# 0.00fF
C4376 sky130_fd_sc_hd__o311a_1_0/A3 sky130_fd_sc_hd__inv_1_49/A 0.09fF
C4377 sky130_fd_sc_hd__dfrtn_1_19/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_761_289# -0.00fF
C4378 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# sky130_fd_sc_hd__inv_1_40/A 0.02fF
C4379 sky130_fd_sc_hd__dfrtn_1_30/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4380 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_37/a_761_289# 0.00fF
C4381 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_37/a_27_47# 0.00fF
C4382 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_37/a_543_47# 0.01fF
C4383 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_37/a_193_47# 0.01fF
C4384 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# DOUT[2] 0.00fF
C4385 sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C4386 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__inv_1_48/A 0.29fF
C4387 sky130_fd_sc_hd__dfrtn_1_8/a_1270_413# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C4388 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__nor3_2_0/A 0.01fF
C4389 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C4390 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_761_289# 0.00fF
C4391 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_543_47# 0.00fF
C4392 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C4393 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_35/a_1108_47# 0.00fF
C4394 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.00fF
C4395 sky130_fd_sc_hd__inv_1_25/A RESET_COUNTERn 0.06fF
C4396 sky130_fd_sc_hd__or2_2_0/X DOUT[23] 0.00fF
C4397 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C4398 sky130_fd_sc_hd__o211a_1_1/a_297_297# DOUT[23] 0.00fF
C4399 DOUT[9] sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.00fF
C4400 sky130_fd_sc_hd__dfrtn_1_38/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C4401 sky130_fd_sc_hd__dfrtn_1_27/a_1270_413# VDD 0.00fF
C4402 sky130_fd_sc_hd__dfrtn_1_27/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4403 sky130_fd_sc_hd__dfrtp_1_3/a_761_289# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.01fF
C4404 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__or2_2_0/a_121_297# 0.00fF
C4405 sky130_fd_sc_hd__nor3_1_18/a_193_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4406 DOUT[1] sky130_fd_sc_hd__dfrtn_1_22/a_193_47# 0.00fF
C4407 sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# RESET_COUNTERn 0.00fF
C4408 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__dfrtn_1_1/a_448_47# 0.00fF
C4409 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__dfrtn_1_1/a_651_413# 0.00fF
C4410 DOUT[2] sky130_fd_sc_hd__inv_1_32/Y 0.01fF
C4411 sky130_fd_sc_hd__dfrtn_1_36/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_651_413# -0.00fF
C4412 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# DOUT[14] 0.01fF
C4413 sky130_fd_sc_hd__o2111a_2_0/a_566_47# RESET_COUNTERn 0.00fF
C4414 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_27_47# 0.01fF
C4415 sky130_fd_sc_hd__inv_1_47/A SEL_CONV_TIME[0] 0.44fF
C4416 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C4417 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C4418 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C4419 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C4420 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C4421 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# VDD 0.15fF
C4422 sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C4423 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_27_47# 0.00fF
C4424 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_193_47# 0.00fF
C4425 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# SEL_CONV_TIME[3] 0.00fF
C4426 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4427 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__nand2_1_1/a_113_47# 0.00fF
C4428 sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C4429 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# VDD 0.00fF
C4430 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_5/a_639_47# 0.00fF
C4431 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.00fF
C4432 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C4433 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C4434 sky130_fd_sc_hd__dfrtn_1_0/a_761_289# sky130_fd_sc_hd__nor3_1_0/A 0.01fF
C4435 sky130_fd_sc_hd__inv_1_7/Y DOUT[19] 0.02fF
C4436 sky130_fd_sc_hd__dfrtp_1_3/a_805_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C4437 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C4438 sky130_fd_sc_hd__dfrtn_1_34/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C4439 sky130_fd_sc_hd__dfrtn_1_12/a_1217_47# VDD 0.00fF
C4440 sky130_fd_sc_hd__dfrtn_1_12/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4441 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C4442 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_30/a_639_47# 0.00fF
C4443 sky130_fd_sc_hd__nor3_2_2/A sky130_fd_sc_hd__inv_1_40/Y 0.05fF
C4444 sky130_fd_sc_hd__dfrtn_1_28/a_193_47# RESET_COUNTERn -0.02fF
C4445 sky130_fd_sc_hd__dfrtn_1_28/a_448_47# DOUT[21] 0.01fF
C4446 sky130_fd_sc_hd__dfrtn_1_33/a_805_47# DOUT[23] 0.00fF
C4447 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# sky130_fd_sc_hd__nor3_1_1/a_109_297# 0.00fF
C4448 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# sky130_fd_sc_hd__nor3_1_1/a_193_297# 0.00fF
C4449 sky130_fd_sc_hd__dfrtn_1_39/a_761_289# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C4450 sky130_fd_sc_hd__dfrtn_1_30/a_761_289# sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C4451 sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# RESET_COUNTERn 0.00fF
C4452 sky130_fd_sc_hd__mux4_1_0/a_750_97# SEL_CONV_TIME[0] 0.03fF
C4453 sky130_fd_sc_hd__dfrtn_1_42/a_805_47# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C4454 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_34/a_1217_47# 0.00fF
C4455 sky130_fd_sc_hd__or3b_2_0/a_472_297# SEL_CONV_TIME[1] 0.00fF
C4456 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_4/Y 0.03fF
C4457 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# DOUT[2] 0.00fF
C4458 sky130_fd_sc_hd__inv_1_14/A sky130_fd_sc_hd__inv_1_0/Y 0.01fF
C4459 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# SEL_CONV_TIME[2] 0.03fF
C4460 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# VIN 0.00fF
C4461 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__or3b_2_0/a_27_47# -0.00fF
C4462 sky130_fd_sc_hd__dfrtn_1_32/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.00fF
C4463 sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C4464 sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# sky130_fd_sc_hd__inv_1_40/A 0.00fF
C4465 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__inv_1_3/Y 0.16fF
C4466 sky130_fd_sc_hd__dfrtn_1_14/a_651_413# DOUT[22] 0.00fF
C4467 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C4468 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C4469 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C4470 sky130_fd_sc_hd__dfrtn_1_32/a_27_47# sky130_fd_sc_hd__inv_1_9/A 0.05fF
C4471 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C4472 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_37/a_651_413# 0.00fF
C4473 sky130_fd_sc_hd__dfrtn_1_24/a_1462_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C4474 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__dfrtn_1_34/a_448_47# 0.00fF
C4475 DOUT[1] sky130_fd_sc_hd__dfrtn_1_23/a_761_289# 0.00fF
C4476 sky130_fd_sc_hd__dfrtn_1_18/a_27_47# DOUT[2] 0.03fF
C4477 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__nor3_2_3/C 0.04fF
C4478 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__nor3_2_0/A 0.03fF
C4479 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# VDD 0.02fF
C4480 sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C4481 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__dfrtn_1_2/a_651_413# 0.00fF
C4482 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__dfrtn_1_2/a_639_47# 0.00fF
C4483 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# 0.00fF
C4484 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# 0.00fF
C4485 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# sky130_fd_sc_hd__dfrtn_1_2/a_543_47# 0.00fF
C4486 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# 0.00fF
C4487 sky130_fd_sc_hd__dfrtn_1_22/a_448_47# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C4488 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_24/a_639_47# -0.00fF
C4489 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_24/a_805_47# -0.00fF
C4490 sky130_fd_sc_hd__o2111a_2_0/a_386_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4491 sky130_fd_sc_hd__o221ai_1_0/a_493_297# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C4492 sky130_fd_sc_hd__nor3_1_12/a_193_297# VDD 0.00fF
C4493 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C4494 sky130_fd_sc_hd__dfrtn_1_39/a_805_47# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C4495 sky130_fd_sc_hd__or3b_2_0/a_388_297# VDD 0.00fF
C4496 DOUT[1] sky130_fd_sc_hd__dfrtn_1_22/a_1462_47# 0.00fF
C4497 sky130_fd_sc_hd__dfrtn_1_31/a_543_47# SEL_CONV_TIME[1] 0.00fF
C4498 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# -0.00fF
C4499 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# 0.00fF
C4500 sky130_fd_sc_hd__mux4_1_0/a_27_413# RESET_COUNTERn 0.01fF
C4501 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4502 DOUT[4] sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C4503 sky130_fd_sc_hd__dfrtn_1_10/a_1283_21# RESET_COUNTERn 0.00fF
C4504 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_41/a_1270_413# 0.00fF
C4505 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_19/a_1108_47# 0.01fF
C4506 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_31/a_193_47# 0.00fF
C4507 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_27_47# 0.00fF
C4508 sky130_fd_sc_hd__dfrtn_1_26/a_805_47# DOUT[23] 0.00fF
C4509 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# DOUT[14] 0.00fF
C4510 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# DOUT[19] 0.00fF
C4511 sky130_fd_sc_hd__inv_1_21/Y DOUT[10] 0.00fF
C4512 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__dfrtn_1_15/a_761_289# 0.00fF
C4513 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_805_47# 0.00fF
C4514 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# 0.00fF
C4515 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# 0.00fF
C4516 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C4517 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# 0.00fF
C4518 sky130_fd_sc_hd__dfrtn_1_25/a_639_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C4519 sky130_fd_sc_hd__dfrtn_1_17/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4520 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C4521 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_805_47# 0.00fF
C4522 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# 0.00fF
C4523 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# 0.00fF
C4524 sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C4525 sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# VDD 0.10fF
C4526 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C4527 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__inv_1_8/A 0.01fF
C4528 sky130_fd_sc_hd__inv_1_26/A outb 0.02fF
C4529 sky130_fd_sc_hd__dfrtn_1_14/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4530 sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# VDD 0.00fF
C4531 sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# DOUT[2] 0.01fF
C4532 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__inv_1_31/A 0.00fF
C4533 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_21/a_1462_47# 0.00fF
C4534 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# 0.00fF
C4535 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# 0.00fF
C4536 sky130_fd_sc_hd__dfrtn_1_12/a_651_413# sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# 0.00fF
C4537 sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# SEL_CONV_TIME[3] 0.00fF
C4538 sky130_fd_sc_hd__nor3_1_4/a_109_297# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C4539 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__o2111a_2_0/a_386_47# 0.00fF
C4540 sky130_fd_sc_hd__or3_1_0/a_183_297# sky130_fd_sc_hd__o2111a_2_0/a_80_21# 0.00fF
C4541 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__o2111a_2_0/a_80_21# 0.00fF
C4542 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__o2111a_2_0/a_386_47# 0.00fF
C4543 sky130_fd_sc_hd__inv_1_29/A CLK_REF 0.01fF
C4544 sky130_fd_sc_hd__nor3_2_3/a_27_297# sky130_fd_sc_hd__dfrtn_1_42/a_448_47# 0.00fF
C4545 sky130_fd_sc_hd__inv_1_45/A SEL_CONV_TIME[1] 0.01fF
C4546 sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C4547 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__dfrtp_1_1/D -0.00fF
C4548 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__inv_1_5/A 0.00fF
C4549 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__inv_1_37/A 0.03fF
C4550 sky130_fd_sc_hd__inv_1_13/Y sky130_fd_sc_hd__inv_1_12/A 0.02fF
C4551 sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C4552 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C4553 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.02fF
C4554 sky130_fd_sc_hd__o311a_1_0/a_266_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C4555 sky130_fd_sc_hd__o211a_1_1/a_215_47# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C4556 sky130_fd_sc_hd__o211a_1_0/a_297_297# DOUT[15] 0.00fF
C4557 sky130_fd_sc_hd__o311a_1_0/a_266_297# SEL_CONV_TIME[0] 0.00fF
C4558 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__nand3b_1_1/a_53_93# 0.00fF
C4559 sky130_fd_sc_hd__dfrtn_1_28/a_1462_47# RESET_COUNTERn 0.00fF
C4560 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C4561 sky130_fd_sc_hd__dfrtn_1_31/a_761_289# VDD 0.06fF
C4562 sky130_fd_sc_hd__inv_1_9/Y DOUT[12] 0.01fF
C4563 sky130_fd_sc_hd__dfrtn_1_0/a_761_289# sky130_fd_sc_hd__nor3_1_1/a_109_297# 0.00fF
C4564 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__nand3b_1_1/Y 0.01fF
C4565 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# sky130_fd_sc_hd__nor3_1_1/a_193_297# 0.00fF
C4566 sky130_fd_sc_hd__mux4_2_0/a_288_47# SEL_CONV_TIME[0] 0.01fF
C4567 sky130_fd_sc_hd__dfrtn_1_35/a_193_47# RESET_COUNTERn -0.02fF
C4568 sky130_fd_sc_hd__dfrtn_1_35/a_448_47# DOUT[21] 0.00fF
C4569 sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# RESET_COUNTERn 0.01fF
C4570 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C4571 sky130_fd_sc_hd__inv_1_3/Y VIN 0.02fF
C4572 DOUT[19] DOUT[10] 0.00fF
C4573 sky130_fd_sc_hd__dfrtn_1_3/a_639_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C4574 DOUT[5] DOUT[17] 0.03fF
C4575 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_193_47# -0.15fF
C4576 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# sky130_fd_sc_hd__or2b_1_0/X 0.01fF
C4577 sky130_fd_sc_hd__or2b_1_0/a_219_297# SEL_CONV_TIME[1] 0.01fF
C4578 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C4579 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__inv_1_53/A 0.01fF
C4580 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_651_413# 0.00fF
C4581 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_39/a_761_289# 0.00fF
C4582 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# 0.00fF
C4583 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_1270_413# 0.00fF
C4584 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# 0.00fF
C4585 sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# SEL_CONV_TIME[2] 0.00fF
C4586 sky130_fd_sc_hd__nor3_1_4/a_109_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4587 sky130_fd_sc_hd__dfrtn_1_32/a_1217_47# sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.00fF
C4588 sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# 0.00fF
C4589 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C4590 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__inv_1_5/A 0.01fF
C4591 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C4592 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_19/a_543_47# 0.00fF
C4593 sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# DOUT[22] 0.00fF
C4594 sky130_fd_sc_hd__inv_1_33/A sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C4595 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__inv_1_31/A 0.01fF
C4596 sky130_fd_sc_hd__dfrtn_1_32/a_1217_47# sky130_fd_sc_hd__inv_1_9/A 0.00fF
C4597 sky130_fd_sc_hd__dfrtn_1_20/a_805_47# RESET_COUNTERn 0.00fF
C4598 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.01fF
C4599 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C4600 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__o221ai_1_0/a_493_297# 0.00fF
C4601 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C4602 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# sky130_fd_sc_hd__o221ai_1_0/a_295_297# 0.00fF
C4603 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# sky130_fd_sc_hd__inv_1_29/Y 0.00fF
C4604 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.00fF
C4605 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_18/a_761_289# 0.00fF
C4606 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_651_413# 0.00fF
C4607 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C4608 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# 0.00fF
C4609 sky130_fd_sc_hd__dfrtn_1_18/a_1217_47# DOUT[2] 0.00fF
C4610 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_1270_413# 0.00fF
C4611 sky130_fd_sc_hd__o2111a_2_0/a_566_47# SEL_CONV_TIME[2] 0.00fF
C4612 sky130_fd_sc_hd__dfrtn_1_42/a_1108_47# sky130_fd_sc_hd__inv_1_25/A 0.00fF
C4613 sky130_fd_sc_hd__dfrtn_1_32/a_651_413# VDD 0.01fF
C4614 sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4615 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4616 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C4617 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__inv_1_33/A 0.11fF
C4618 sky130_fd_sc_hd__nor3_2_1/a_27_297# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C4619 outb en 0.00fF
C4620 sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# DOUT[11] 0.00fF
C4621 sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C4622 sky130_fd_sc_hd__dfrtn_1_36/a_448_47# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C4623 CLK_REF DOUT[23] 0.00fF
C4624 sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# sky130_fd_sc_hd__inv_1_52/Y 0.02fF
C4625 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C4626 sky130_fd_sc_hd__dfrtp_1_3/a_543_47# sky130_fd_sc_hd__or2_2_0/A 0.01fF
C4627 sky130_fd_sc_hd__o311a_1_0/a_81_21# DOUT[21] 0.00fF
C4628 sky130_fd_sc_hd__mux4_1_0/a_668_97# RESET_COUNTERn 0.00fF
C4629 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_26/a_448_47# 0.00fF
C4630 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# sky130_fd_sc_hd__inv_1_37/A 0.01fF
C4631 sky130_fd_sc_hd__o2111a_2_0/a_386_47# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C4632 sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# sky130_fd_sc_hd__dfrtn_1_28/a_27_47# 0.01fF
C4633 sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# sky130_fd_sc_hd__dfrtn_1_28/a_193_47# 0.01fF
C4634 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_24/a_448_47# 0.00fF
C4635 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.02fF
C4636 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C4637 sky130_fd_sc_hd__nor3_1_12/a_109_297# sky130_fd_sc_hd__inv_1_9/Y 0.00fF
C4638 sky130_fd_sc_hd__dfrtn_1_34/a_651_413# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C4639 sky130_fd_sc_hd__nor3_2_1/A lc_out 0.07fF
C4640 sky130_fd_sc_hd__dfrtn_1_42/a_543_47# sky130_fd_sc_hd__nor3_2_3/A 0.01fF
C4641 sky130_fd_sc_hd__o211a_1_0/a_215_47# lc_out 0.01fF
C4642 sky130_fd_sc_hd__dfrtn_1_28/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4643 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# DOUT[11] 0.00fF
C4644 sky130_fd_sc_hd__dfrtn_1_0/a_651_413# sky130_fd_sc_hd__nor3_1_0/a_109_297# 0.00fF
C4645 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C4646 sky130_fd_sc_hd__dfrtn_1_0/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4647 sky130_fd_sc_hd__dfrtn_1_14/a_761_289# DOUT[9] 0.00fF
C4648 DOUT[4] sky130_fd_sc_hd__or3b_2_0/X 0.01fF
C4649 sky130_fd_sc_hd__dfrtn_1_32/a_193_47# sky130_fd_sc_hd__dfrtn_1_32/a_805_47# -0.00fF
C4650 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# VDD 0.08fF
C4651 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__inv_1_33/A 0.02fF
C4652 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# RESET_COUNTERn 0.03fF
C4653 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_34/a_193_47# 0.00fF
C4654 sky130_fd_sc_hd__dfrtn_1_22/a_1217_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C4655 sky130_fd_sc_hd__o311a_1_0/a_81_21# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C4656 DOUT[4] sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# 0.00fF
C4657 sky130_fd_sc_hd__nand3b_1_0/a_316_47# DOUT[21] 0.00fF
C4658 sky130_fd_sc_hd__o221ai_1_0/a_295_297# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C4659 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_805_47# 0.00fF
C4660 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# 0.00fF
C4661 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C4662 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C4663 sky130_fd_sc_hd__nor3_1_5/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4664 sky130_fd_sc_hd__dfrtn_1_19/a_761_289# sky130_fd_sc_hd__inv_1_28/A 0.02fF
C4665 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__inv_1_8/Y 0.02fF
C4666 sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# sky130_fd_sc_hd__nor3_1_5/a_193_297# 0.00fF
C4667 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C4668 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C4669 sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C4670 sky130_fd_sc_hd__inv_1_26/A sky130_fd_sc_hd__nor3_2_3/A 0.01fF
C4671 sky130_fd_sc_hd__or2_2_0/B lc_out 0.05fF
C4672 sky130_fd_sc_hd__inv_1_9/Y sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C4673 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C4674 sky130_fd_sc_hd__dfrtn_1_35/a_1462_47# RESET_COUNTERn -0.00fF
C4675 sky130_fd_sc_hd__dfrtn_1_32/a_193_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C4676 sky130_fd_sc_hd__nor3_1_11/a_193_297# RESET_COUNTERn 0.00fF
C4677 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_1/a_193_47# 0.00fF
C4678 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# DOUT[3] 0.00fF
C4679 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_39/a_1462_47# 0.00fF
C4680 sky130_fd_sc_hd__nor3_1_8/a_193_297# VIN 0.00fF
C4681 sky130_fd_sc_hd__dfrtp_1_1/a_639_47# RESET_COUNTERn 0.00fF
C4682 sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__dfrtn_1_25/a_27_47# 0.00fF
C4683 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_25/a_193_47# 0.00fF
C4684 sky130_fd_sc_hd__o2111a_2_0/a_458_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C4685 sky130_fd_sc_hd__dfrtp_1_3/a_651_413# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C4686 sky130_fd_sc_hd__dfrtp_1_3/a_543_47# sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# 0.00fF
C4687 sky130_fd_sc_hd__dfrtp_1_3/a_1283_21# sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# 0.00fF
C4688 sky130_fd_sc_hd__dfrtp_1_3/a_448_47# sky130_fd_sc_hd__dfrtn_1_17/a_761_289# 0.00fF
C4689 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_651_413# 0.00fF
C4690 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C4691 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtp_1_2/a_761_289# -0.00fF
C4692 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__nor3_1_0/A 0.01fF
C4693 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_3/Y 0.02fF
C4694 sky130_fd_sc_hd__dfrtn_1_34/a_1217_47# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C4695 sky130_fd_sc_hd__dfrtn_1_34/a_805_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C4696 DOUT[1] sky130_fd_sc_hd__nor3_2_3/B 0.07fF
C4697 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C4698 sky130_fd_sc_hd__nand3b_1_0/a_316_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C4699 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_7/A 0.01fF
C4700 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4701 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__dfrtn_1_29/a_448_47# 0.00fF
C4702 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# 0.00fF
C4703 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__dfrtn_1_29/a_651_413# 0.00fF
C4704 sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__nor3_2_3/B 0.31fF
C4705 sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# sky130_fd_sc_hd__inv_1_7/A 0.01fF
C4706 sky130_fd_sc_hd__o211a_1_0/a_215_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C4707 sky130_fd_sc_hd__dfrtp_1_3/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4708 sky130_fd_sc_hd__dfrtp_1_3/a_651_413# VDD 0.01fF
C4709 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__nor3_1_12/a_193_297# 0.00fF
C4710 sky130_fd_sc_hd__inv_1_31/Y DOUT[2] 0.00fF
C4711 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_1/a_805_47# -0.00fF
C4712 sky130_fd_sc_hd__dfrtn_1_29/a_639_47# SEL_CONV_TIME[1] 0.00fF
C4713 sky130_fd_sc_hd__dfrtn_1_20/a_543_47# sky130_fd_sc_hd__dfrtn_1_21/a_193_47# 0.00fF
C4714 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C4715 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__inv_1_48/A 0.25fF
C4716 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__dfrtn_1_24/a_27_47# 0.00fF
C4717 sky130_fd_sc_hd__or3b_2_0/a_388_297# sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# 0.00fF
C4718 sky130_fd_sc_hd__or3_1_0/C DOUT[21] 0.01fF
C4719 DOUT[4] sky130_fd_sc_hd__dfrtn_1_34/a_193_47# 0.01fF
C4720 sky130_fd_sc_hd__mux4_2_0/a_1281_47# DOUT[21] 0.00fF
C4721 sky130_fd_sc_hd__mux4_2_0/a_872_316# RESET_COUNTERn 0.00fF
C4722 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__dfrtp_1_1/D 0.00fF
C4723 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__o211a_1_1/a_297_297# 0.00fF
C4724 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# 0.00fF
C4725 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# -0.00fF
C4726 sky130_fd_sc_hd__or2_2_0/B sky130_fd_sc_hd__nor3_2_3/B 0.21fF
C4727 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# -0.00fF
C4728 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__dfrtn_1_13/a_543_47# -0.00fF
C4729 sky130_fd_sc_hd__or2b_1_0/X DOUT[21] 0.01fF
C4730 sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# DOUT[11] 0.00fF
C4731 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# RESET_COUNTERn 0.01fF
C4732 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_10/a_193_47# 0.01fF
C4733 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# DOUT[23] 0.00fF
C4734 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# DOUT[19] 0.00fF
C4735 sky130_fd_sc_hd__dfrtn_1_35/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4736 sky130_fd_sc_hd__nor3_1_15/a_109_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4737 sky130_fd_sc_hd__dfrtn_1_8/a_193_47# DOUT[12] 0.00fF
C4738 sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# RESET_COUNTERn 0.00fF
C4739 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_34/a_1462_47# 0.00fF
C4740 sky130_fd_sc_hd__dfrtp_1_3/a_448_47# sky130_fd_sc_hd__nor3_2_1/a_27_297# 0.00fF
C4741 sky130_fd_sc_hd__dfrtn_1_18/a_193_47# sky130_fd_sc_hd__inv_1_27/Y 0.00fF
C4742 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C4743 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__inv_1_53/A 0.02fF
C4744 sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# VDD 0.00fF
C4745 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C4746 sky130_fd_sc_hd__o311a_1_0/A3 sky130_fd_sc_hd__or3_1_0/C 0.00fF
C4747 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C4748 sky130_fd_sc_hd__mux4_2_0/a_1281_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C4749 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4750 CLK_REF sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.01fF
C4751 sky130_fd_sc_hd__nor3_2_3/a_281_297# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C4752 sky130_fd_sc_hd__dfrtn_1_3/a_1462_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C4753 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__o211a_1_1/a_297_297# 0.00fF
C4754 DOUT[9] sky130_fd_sc_hd__inv_1_7/A 0.02fF
C4755 sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# sky130_fd_sc_hd__dfrtn_1_18/a_543_47# 0.00fF
C4756 sky130_fd_sc_hd__dfrtn_1_20/a_651_413# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C4757 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_448_47# 0.00fF
C4758 sky130_fd_sc_hd__dfrtn_1_18/a_27_47# sky130_fd_sc_hd__inv_1_30/Y 0.01fF
C4759 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C4760 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__o2111a_2_0/X 0.02fF
C4761 sky130_fd_sc_hd__nor3_1_1/a_193_297# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C4762 sky130_fd_sc_hd__dfrtn_1_32/a_1462_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C4763 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_34/a_193_47# 0.00fF
C4764 sky130_fd_sc_hd__or2b_1_0/X sky130_fd_sc_hd__o311a_1_0/A3 0.04fF
C4765 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__o211a_1_0/a_79_21# 0.01fF
C4766 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__inv_1_11/A 0.12fF
C4767 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_448_47# 0.00fF
C4768 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# sky130_fd_sc_hd__dfrtn_1_36/a_543_47# 0.00fF
C4769 sky130_fd_sc_hd__dfrtn_1_23/a_651_413# sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C4770 sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# sky130_fd_sc_hd__dfrtn_1_36/a_761_289# 0.00fF
C4771 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_651_413# 0.00fF
C4772 sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# RESET_COUNTERn 0.04fF
C4773 sky130_fd_sc_hd__dfrtn_1_27/a_639_47# DOUT[21] 0.00fF
C4774 sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C4775 sky130_fd_sc_hd__dfrtn_1_19/a_1462_47# sky130_fd_sc_hd__inv_1_35/Y 0.00fF
C4776 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C4777 sky130_fd_sc_hd__dfrtn_1_35/a_1108_47# sky130_fd_sc_hd__inv_1_38/A 0.01fF
C4778 sky130_fd_sc_hd__dfrtn_1_3/a_805_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C4779 sky130_fd_sc_hd__dfrtn_1_11/a_1270_413# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C4780 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C4781 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__dfrtn_1_25/a_651_413# 0.00fF
C4782 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_25/a_639_47# 0.00fF
C4783 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_32/a_651_413# 0.00fF
C4784 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C4785 sky130_fd_sc_hd__dfrtn_1_30/a_761_289# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C4786 sky130_fd_sc_hd__nor3_2_0/a_281_297# sky130_fd_sc_hd__dfrtn_1_12/a_193_47# 0.00fF
C4787 sky130_fd_sc_hd__o311a_1_0/a_585_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4788 DOUT[13] sky130_fd_sc_hd__dfrtn_1_30/a_27_47# 0.02fF
C4789 sky130_fd_sc_hd__dfrtn_1_37/a_805_47# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C4790 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# sky130_fd_sc_hd__mux4_2_0/a_600_345# 0.00fF
C4791 sky130_fd_sc_hd__dfrtn_1_37/a_1270_413# sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.00fF
C4792 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# sky130_fd_sc_hd__mux4_2_0/a_193_47# 0.00fF
C4793 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C4794 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# sky130_fd_sc_hd__mux4_2_0/a_372_413# 0.00fF
C4795 sky130_fd_sc_hd__dfrtn_1_38/a_543_47# DOUT[2] 0.00fF
C4796 sky130_fd_sc_hd__dfrtn_1_4/a_1270_413# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C4797 sky130_fd_sc_hd__mux4_2_0/a_600_345# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4798 sky130_fd_sc_hd__dfrtn_1_42/a_193_47# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C4799 sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__inv_1_22/A 0.00fF
C4800 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C4801 sky130_fd_sc_hd__inv_1_0/A DOUT[4] 0.00fF
C4802 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_0/Y 0.14fF
C4803 sky130_fd_sc_hd__dfrtn_1_10/a_1270_413# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C4804 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__inv_1_32/A 0.20fF
C4805 sky130_fd_sc_hd__dfrtn_1_36/a_193_47# DOUT[21] 0.02fF
C4806 sky130_fd_sc_hd__dfrtn_1_29/a_805_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C4807 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__dfrtn_1_24/a_1270_413# 0.00fF
C4808 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__dfrtn_1_24/a_1462_47# 0.00fF
C4809 sky130_fd_sc_hd__dfrtn_1_21/a_1217_47# VDD 0.00fF
C4810 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# RESET_COUNTERn 0.01fF
C4811 sky130_fd_sc_hd__dfrtn_1_9/a_543_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C4812 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# 0.00fF
C4813 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# sky130_fd_sc_hd__inv_1_0/Y 0.01fF
C4814 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C4815 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__nor3_1_1/a_109_297# 0.00fF
C4816 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# VDD 0.09fF
C4817 sky130_fd_sc_hd__dfrtn_1_4/a_448_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C4818 sky130_fd_sc_hd__inv_1_25/A sky130_fd_sc_hd__nor3_2_2/A 0.03fF
C4819 sky130_fd_sc_hd__dfrtn_1_22/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4820 sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4821 sky130_fd_sc_hd__dfrtn_1_12/a_651_413# RESET_COUNTERn 0.00fF
C4822 sky130_fd_sc_hd__dfrtn_1_39/a_543_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C4823 sky130_fd_sc_hd__dfrtn_1_38/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# -0.00fF
C4824 sky130_fd_sc_hd__dfrtn_1_38/a_761_289# sky130_fd_sc_hd__dfrtn_1_38/a_543_47# -0.00fF
C4825 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# -0.00fF
C4826 sky130_fd_sc_hd__dfrtn_1_20/a_651_413# sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# 0.00fF
C4827 sky130_fd_sc_hd__dfrtn_1_22/a_639_47# VDD 0.00fF
C4828 DOUT[1] sky130_fd_sc_hd__dfrtn_1_42/a_651_413# 0.00fF
C4829 sky130_fd_sc_hd__nor3_1_12/a_109_297# sky130_fd_sc_hd__dfrtn_1_8/a_193_47# 0.00fF
C4830 sky130_fd_sc_hd__nor3_1_12/a_193_297# sky130_fd_sc_hd__dfrtn_1_8/a_27_47# 0.00fF
C4831 sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C4832 sky130_fd_sc_hd__dfrtn_1_28/a_1217_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C4833 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__dfrtn_1_21/a_651_413# -0.00fF
C4834 sky130_fd_sc_hd__dfrtn_1_21/a_448_47# sky130_fd_sc_hd__dfrtn_1_21/a_193_47# -0.00fF
C4835 outb VIN 1.36fF
C4836 DOUT[4] sky130_fd_sc_hd__dfrtn_1_34/a_1462_47# 0.00fF
C4837 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__dfrtn_1_25/a_193_47# 0.00fF
C4838 sky130_fd_sc_hd__nand3b_1_0/a_232_47# sky130_fd_sc_hd__dfrtn_1_25/a_27_47# 0.00fF
C4839 DOUT[19] sky130_fd_sc_hd__inv_1_4/Y 0.05fF
C4840 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C4841 sky130_fd_sc_hd__dfrtn_1_18/a_543_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C4842 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__dfrtn_1_6/a_448_47# 0.00fF
C4843 sky130_fd_sc_hd__nor3_1_11/a_109_297# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C4844 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C4845 sky130_fd_sc_hd__dfrtn_1_23/a_805_47# sky130_fd_sc_hd__inv_1_40/A 0.00fF
C4846 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# 0.00fF
C4847 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# sky130_fd_sc_hd__dfrtp_1_1/a_761_289# 0.00fF
C4848 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# 0.00fF
C4849 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# 0.01fF
C4850 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__mux4_2_0/a_600_345# 0.00fF
C4851 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C4852 sky130_fd_sc_hd__o211a_1_1/a_215_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C4853 sky130_fd_sc_hd__nor3_1_5/A DOUT[22] 0.02fF
C4854 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_26/a_543_47# 0.00fF
C4855 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__inv_1_1/A 0.09fF
C4856 sky130_fd_sc_hd__dfrtn_1_8/a_651_413# sky130_fd_sc_hd__inv_1_9/A 0.00fF
C4857 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_10/a_1462_47# 0.00fF
C4858 sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# DOUT[23] 0.00fF
C4859 sky130_fd_sc_hd__dfrtn_1_26/a_448_47# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C4860 sky130_fd_sc_hd__dfrtn_1_26/a_543_47# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C4861 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_651_413# 0.00fF
C4862 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__inv_1_5/A 0.01fF
C4863 sky130_fd_sc_hd__dfrtn_1_8/a_1462_47# DOUT[12] 0.00fF
C4864 sky130_fd_sc_hd__dfrtn_1_3/a_639_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C4865 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C4866 sky130_fd_sc_hd__mux4_2_0/a_872_316# SEL_CONV_TIME[3] 0.01fF
C4867 sky130_fd_sc_hd__dfrtn_1_16/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C4868 sky130_fd_sc_hd__dfrtn_1_27/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C4869 sky130_fd_sc_hd__dfrtn_1_16/a_651_413# VDD 0.01fF
C4870 sky130_fd_sc_hd__dfrtn_1_8/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.13fF
C4871 sky130_fd_sc_hd__dfrtn_1_8/a_543_47# VDD 0.05fF
C4872 sky130_fd_sc_hd__nor3_1_3/a_109_297# DOUT[14] 0.00fF
C4873 sky130_fd_sc_hd__dfrtn_1_18/a_1462_47# sky130_fd_sc_hd__inv_1_27/Y 0.00fF
C4874 sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C4875 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_761_289# -0.00fF
C4876 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_805_47# -0.00fF
C4877 sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C4878 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# sky130_fd_sc_hd__inv_1_47/A 0.01fF
C4879 CLK_REF sky130_fd_sc_hd__dfrtn_1_19/a_1462_47# 0.00fF
C4880 DOUT[23] sky130_fd_sc_hd__inv_1_43/A 0.00fF
C4881 sky130_fd_sc_hd__dfrtn_1_21/a_193_47# sky130_fd_sc_hd__inv_1_35/A 0.01fF
C4882 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C4883 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# 0.01fF
C4884 sky130_fd_sc_hd__dfrtn_1_18/a_1217_47# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C4885 sky130_fd_sc_hd__nor3_1_13/a_109_297# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C4886 sky130_fd_sc_hd__dfrtn_1_31/a_1283_21# SEL_CONV_TIME[0] 0.01fF
C4887 SEL_CONV_TIME[1] RESET_COUNTERn 0.38fF
C4888 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C4889 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# DOUT[2] 0.00fF
C4890 sky130_fd_sc_hd__dfrtp_1_0/a_639_47# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C4891 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C4892 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_40/a_448_47# -0.00fF
C4893 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# -0.00fF
C4894 sky130_fd_sc_hd__inv_1_3/A DOUT[6] 0.17fF
C4895 sky130_fd_sc_hd__nor3_2_1/A DOUT[0] 0.00fF
C4896 sky130_fd_sc_hd__dfrtn_1_23/a_1462_47# sky130_fd_sc_hd__dfrtn_1_36/a_448_47# 0.00fF
C4897 sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C4898 sky130_fd_sc_hd__o211a_1_0/a_215_47# DOUT[0] 0.00fF
C4899 sky130_fd_sc_hd__o211a_1_0/a_510_47# out 0.00fF
C4900 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__inv_1_13/Y 0.13fF
C4901 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4902 sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C4903 sky130_fd_sc_hd__nor3_1_11/a_193_297# HEADER_0/a_508_138# 0.00fF
C4904 sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# sky130_fd_sc_hd__inv_1_8/Y 0.01fF
C4905 sky130_fd_sc_hd__mux4_2_0/a_872_316# SEL_CONV_TIME[2] 0.00fF
C4906 sky130_fd_sc_hd__nor3_1_11/a_193_297# sky130_fd_sc_hd__dfrtn_1_2/a_448_47# 0.00fF
C4907 sky130_fd_sc_hd__dfrtn_1_23/a_805_47# VDD 0.00fF
C4908 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4909 DOUT[13] sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# 0.00fF
C4910 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# 0.00fF
C4911 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_805_47# 0.00fF
C4912 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C4913 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__dfrtn_1_38/a_761_289# 0.00fF
C4914 DOUT[9] sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C4915 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_3/a_543_47# 0.00fF
C4916 sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4917 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__or3b_2_0/a_176_21# 0.00fF
C4918 sky130_fd_sc_hd__dfrtn_1_7/a_448_47# VDD 0.01fF
C4919 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# RESET_COUNTERn 0.02fF
C4920 sky130_fd_sc_hd__dfrtn_1_42/a_1462_47# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C4921 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# DOUT[14] 0.00fF
C4922 sky130_fd_sc_hd__dfrtn_1_9/a_761_289# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C4923 sky130_fd_sc_hd__dfrtn_1_36/a_651_413# RESET_COUNTERn 0.00fF
C4924 sky130_fd_sc_hd__dfrtn_1_36/a_1462_47# DOUT[21] 0.00fF
C4925 sky130_fd_sc_hd__dfrtn_1_37/a_1462_47# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C4926 sky130_fd_sc_hd__inv_1_37/A sky130_fd_sc_hd__inv_1_6/A 0.00fF
C4927 sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C4928 DOUT[4] sky130_fd_sc_hd__dfrtn_1_28/a_1108_47# 0.00fF
C4929 sky130_fd_sc_hd__dfrtp_1_0/a_639_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C4930 sky130_fd_sc_hd__or2_2_0/B DOUT[0] 0.00fF
C4931 sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C4932 sky130_fd_sc_hd__o311a_1_0/a_585_47# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C4933 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# VDD 0.00fF
C4934 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4935 sky130_fd_sc_hd__nor3_2_3/C DOUT[6] 0.03fF
C4936 VDD DOUT[8] 0.42fF
C4937 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C4938 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C4939 sky130_fd_sc_hd__mux4_2_0/a_600_345# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C4940 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C4941 sky130_fd_sc_hd__or3b_2_0/a_472_297# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C4942 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C4943 sky130_fd_sc_hd__dfrtn_1_21/a_543_47# sky130_fd_sc_hd__inv_1_35/Y 0.01fF
C4944 sky130_fd_sc_hd__or2b_1_0/a_27_53# SEL_CONV_TIME[0] 0.02fF
C4945 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C4946 sky130_fd_sc_hd__dfrtn_1_40/a_1462_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C4947 sky130_fd_sc_hd__dfrtn_1_27/a_651_413# DOUT[23] 0.00fF
C4948 CLK_REF sky130_fd_sc_hd__or2_2_0/X 0.32fF
C4949 sky130_fd_sc_hd__nor3_1_13/a_109_297# sky130_fd_sc_hd__dfrtn_1_10/a_27_47# 0.00fF
C4950 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# DOUT[0] 0.00fF
C4951 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# 0.00fF
C4952 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C4953 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C4954 CLK_REF sky130_fd_sc_hd__o211a_1_1/a_297_297# 0.00fF
C4955 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C4956 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# SEL_CONV_TIME[1] 0.00fF
C4957 sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# 0.00fF
C4958 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# 0.01fF
C4959 sky130_fd_sc_hd__dfrtn_1_25/a_651_413# sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.00fF
C4960 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_651_413# 0.00fF
C4961 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_1270_413# 0.00fF
C4962 sky130_fd_sc_hd__dfrtn_1_25/a_448_47# sky130_fd_sc_hd__dfrtn_1_27/a_761_289# 0.00fF
C4963 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_31/a_27_47# 0.00fF
C4964 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C4965 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C4966 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__dfrtn_1_13/a_651_413# 0.00fF
C4967 sky130_fd_sc_hd__nor3_1_4/a_193_297# DOUT[6] 0.00fF
C4968 sky130_fd_sc_hd__nor3_1_4/a_109_297# DOUT[7] 0.00fF
C4969 sky130_fd_sc_hd__dfrtn_1_42/a_448_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C4970 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C4971 sky130_fd_sc_hd__dfrtn_1_8/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C4972 sky130_fd_sc_hd__nor3_1_14/a_193_297# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C4973 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C4974 sky130_fd_sc_hd__dfrtn_1_34/a_639_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C4975 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C4976 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C4977 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C4978 sky130_fd_sc_hd__dfrtn_1_32/a_543_47# RESET_COUNTERn 0.00fF
C4979 sky130_fd_sc_hd__dfrtn_1_32/a_1270_413# DOUT[21] 0.00fF
C4980 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__dfrtn_1_33/a_27_47# 0.00fF
C4981 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__dfrtn_1_34/a_448_47# 0.00fF
C4982 sky130_fd_sc_hd__dfrtn_1_31/a_543_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C4983 sky130_fd_sc_hd__dfrtn_1_8/a_761_289# sky130_fd_sc_hd__inv_1_9/Y 0.01fF
C4984 sky130_fd_sc_hd__dfrtn_1_28/a_193_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C4985 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# CLK_REF 0.00fF
C4986 DOUT[4] sky130_fd_sc_hd__dfrtn_1_10/a_1270_413# 0.00fF
C4987 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C4988 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__dfrtn_1_22/a_1283_21# -0.00fF
C4989 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# sky130_fd_sc_hd__dfrtn_1_22/a_543_47# -0.00fF
C4990 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__or3b_2_0/a_27_47# 0.03fF
C4991 sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C4992 sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C4993 sky130_fd_sc_hd__dfrtn_1_24/a_448_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C4994 sky130_fd_sc_hd__or2b_1_0/a_219_297# DOUT[21] 0.00fF
C4995 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# VDD 0.06fF
C4996 VDD sky130_fd_sc_hd__inv_1_43/Y 0.26fF
C4997 sky130_fd_sc_hd__dfrtn_1_25/a_805_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C4998 sky130_fd_sc_hd__nor3_1_0/a_193_297# VDD 0.00fF
C4999 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_17/a_543_47# 0.01fF
C5000 sky130_fd_sc_hd__dfrtn_1_39/a_448_47# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C5001 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# VDD 0.07fF
C5002 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__mux4_2_0/a_397_47# 0.00fF
C5003 SEL_CONV_TIME[1] SEL_CONV_TIME[3] 0.08fF
C5004 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C5005 sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# RESET_COUNTERn 0.00fF
C5006 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__o2111a_2_0/a_458_47# -0.00fF
C5007 sky130_fd_sc_hd__dfrtn_1_41/a_805_47# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C5008 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# RESET_COUNTERn 0.04fF
C5009 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.01fF
C5010 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5011 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__nor3_2_3/C 0.37fF
C5012 sky130_fd_sc_hd__inv_1_17/A sky130_fd_sc_hd__inv_1_23/A 0.18fF
C5013 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C5014 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# sky130_fd_sc_hd__inv_1_38/A 0.00fF
C5015 CLK_REF sky130_fd_sc_hd__dfrtn_1_21/a_543_47# 0.01fF
C5016 sky130_fd_sc_hd__dfrtn_1_19/a_543_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C5017 sky130_fd_sc_hd__dfrtn_1_0/a_639_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C5018 DOUT[4] sky130_fd_sc_hd__dfrtn_1_35/a_1108_47# 0.01fF
C5019 sky130_fd_sc_hd__dfrtn_1_11/a_805_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C5020 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# 0.00fF
C5021 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# 0.00fF
C5022 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# 0.00fF
C5023 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_31/a_193_47# 0.00fF
C5024 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C5025 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C5026 sky130_fd_sc_hd__dfrtn_1_31/a_639_47# RESET_COUNTERn 0.00fF
C5027 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C5028 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.00fF
C5029 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__dfrtn_1_26/a_761_289# 0.00fF
C5030 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C5031 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__dfrtn_1_28/a_27_47# 0.00fF
C5032 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C5033 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# 0.00fF
C5034 sky130_fd_sc_hd__inv_1_15/A sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C5035 SEL_CONV_TIME[1] SEL_CONV_TIME[2] 0.01fF
C5036 sky130_fd_sc_hd__dfrtn_1_9/a_639_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C5037 sky130_fd_sc_hd__dfrtn_1_32/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5038 sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# SEL_CONV_TIME[1] 0.00fF
C5039 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C5040 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# 0.00fF
C5041 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C5042 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_8/a_543_47# 0.01fF
C5043 sky130_fd_sc_hd__dfrtn_1_19/a_27_47# sky130_fd_sc_hd__inv_1_28/Y 0.02fF
C5044 sky130_fd_sc_hd__dfrtn_1_20/a_1270_413# DOUT[2] 0.00fF
C5045 sky130_fd_sc_hd__inv_1_29/Y sky130_fd_sc_hd__inv_1_28/Y 0.01fF
C5046 outb sky130_fd_sc_hd__inv_1_11/A 0.00fF
C5047 sky130_fd_sc_hd__inv_1_19/A en 0.01fF
C5048 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# DOUT[3] 0.02fF
C5049 sky130_fd_sc_hd__dfrtn_1_31/a_651_413# DONE 0.00fF
C5050 sky130_fd_sc_hd__o221ai_1_0/a_295_297# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C5051 sky130_fd_sc_hd__mux4_2_0/a_397_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C5052 sky130_fd_sc_hd__dfrtn_1_9/a_448_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C5053 sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# sky130_fd_sc_hd__inv_1_27/Y 0.00fF
C5054 CLK_REF sky130_fd_sc_hd__inv_1_35/Y 0.06fF
C5055 sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C5056 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__inv_1_2/A 0.08fF
C5057 sky130_fd_sc_hd__dfrtn_1_29/a_805_47# SEL_CONV_TIME[0] 0.00fF
C5058 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_33/a_651_413# 0.00fF
C5059 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__dfrtn_1_33/a_193_47# 0.00fF
C5060 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_33/a_805_47# 0.00fF
C5061 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__dfrtn_1_33/a_1108_47# 0.00fF
C5062 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.00fF
C5063 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__or2_2_0/X 0.01fF
C5064 sky130_fd_sc_hd__dfrtp_1_3/a_543_47# RESET_COUNTERn 0.01fF
C5065 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__inv_1_54/Y 0.02fF
C5066 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__o211a_1_1/a_297_297# 0.00fF
C5067 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.00fF
C5068 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__o211a_1_1/a_215_47# 0.00fF
C5069 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C5070 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C5071 sky130_fd_sc_hd__nor3_2_3/C DOUT[23] 0.78fF
C5072 sky130_fd_sc_hd__dfrtn_1_17/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5073 sky130_fd_sc_hd__dfrtn_1_10/a_1270_413# outb 0.00fF
C5074 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C5075 DOUT[1] DOUT[2] 0.00fF
C5076 sky130_fd_sc_hd__mux4_1_0/a_27_47# DOUT[2] 0.00fF
C5077 sky130_fd_sc_hd__nor3_1_10/a_109_297# DOUT[14] 0.00fF
C5078 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C5079 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# VDD 0.03fF
C5080 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C5081 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__inv_1_53/A 0.02fF
C5082 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_761_289# 0.00fF
C5083 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_3/a_193_47# 0.00fF
C5084 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__dfrtn_1_3/a_27_47# 0.00fF
C5085 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C5086 sky130_fd_sc_hd__dfrtn_1_12/a_639_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C5087 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__inv_1_46/Y 0.00fF
C5088 sky130_fd_sc_hd__dfrtn_1_20/a_761_289# sky130_fd_sc_hd__inv_1_35/Y 0.00fF
C5089 sky130_fd_sc_hd__nor3_1_17/a_109_297# sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# 0.00fF
C5090 sky130_fd_sc_hd__dfrtn_1_3/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5091 sky130_fd_sc_hd__dfrtn_1_3/a_1462_47# VDD 0.00fF
C5092 sky130_fd_sc_hd__dfrtn_1_14/a_805_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C5093 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# 0.00fF
C5094 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# 0.00fF
C5095 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__dfrtp_1_2/a_193_47# 0.00fF
C5096 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_2/a_651_413# 0.00fF
C5097 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# 0.00fF
C5098 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__inv_1_4/A 0.00fF
C5099 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__nor3_2_3/B 0.03fF
C5100 sky130_fd_sc_hd__dfrtn_1_34/a_1270_413# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C5101 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C5102 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C5103 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C5104 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C5105 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C5106 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_805_47# 0.00fF
C5107 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# 0.00fF
C5108 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__inv_1_53/Y 0.06fF
C5109 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# RESET_COUNTERn 0.00fF
C5110 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__inv_1_44/Y 0.53fF
C5111 sky130_fd_sc_hd__dfrtn_1_42/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C5112 sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# VDD 0.08fF
C5113 sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# sky130_fd_sc_hd__inv_1_38/A 0.00fF
C5114 sky130_fd_sc_hd__nand3b_1_1/Y sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C5115 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__nor3_2_0/A 0.01fF
C5116 sky130_fd_sc_hd__nor3_1_16/a_109_297# VDD 0.00fF
C5117 DOUT[4] sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C5118 HEADER_1/a_508_138# sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# 0.00fF
C5119 sky130_fd_sc_hd__dfrtn_1_29/a_639_47# DOUT[21] 0.00fF
C5120 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# RESET_COUNTERn 0.01fF
C5121 sky130_fd_sc_hd__or2_2_0/a_39_297# sky130_fd_sc_hd__o211a_1_1/X 0.00fF
C5122 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C5123 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.03fF
C5124 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.01fF
C5125 sky130_fd_sc_hd__nor3_2_1/a_281_297# DOUT[23] 0.00fF
C5126 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# -0.00fF
C5127 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__dfrtn_1_23/a_448_47# -0.00fF
C5128 sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C5129 sky130_fd_sc_hd__inv_1_0/Y DOUT[17] 0.00fF
C5130 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C5131 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C5132 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# VDD 0.06fF
C5133 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_9/A 0.27fF
C5134 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C5135 sky130_fd_sc_hd__dfrtn_1_4/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5136 sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C5137 sky130_fd_sc_hd__dfrtn_1_4/a_1270_413# VDD 0.00fF
C5138 sky130_fd_sc_hd__dfrtn_1_14/a_448_47# DOUT[11] 0.00fF
C5139 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C5140 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# 0.00fF
C5141 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# 0.00fF
C5142 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_26/a_805_47# 0.00fF
C5143 sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__dfrtn_1_26/a_543_47# 0.00fF
C5144 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__inv_1_31/A 0.00fF
C5145 sky130_fd_sc_hd__dfrtn_1_7/a_448_47# DOUT[3] 0.00fF
C5146 sky130_fd_sc_hd__nor3_1_9/a_109_297# DOUT[14] 0.00fF
C5147 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.01fF
C5148 SLC_0/a_438_293# VDD 0.08fF
C5149 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C5150 sky130_fd_sc_hd__dfrtn_1_19/a_1217_47# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C5151 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# DOUT[15] 0.62fF
C5152 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# sky130_fd_sc_hd__dfrtn_1_16/a_1217_47# -0.00fF
C5153 sky130_fd_sc_hd__dfrtn_1_7/a_448_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C5154 sky130_fd_sc_hd__dfrtn_1_8/a_27_47# sky130_fd_sc_hd__dfrtn_1_8/a_543_47# -0.00fF
C5155 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# DOUT[21] 0.00fF
C5156 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# DOUT[3] 0.00fF
C5157 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__nor3_1_2/a_109_297# 0.00fF
C5158 DOUT[8] DOUT[3] 0.00fF
C5159 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C5160 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.00fF
C5161 sky130_fd_sc_hd__inv_1_6/A DOUT[14] 0.91fF
C5162 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C5163 sky130_fd_sc_hd__dfrtn_1_29/a_639_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C5164 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# sky130_fd_sc_hd__dfrtn_1_7/a_761_289# 0.01fF
C5165 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__dfrtn_1_7/a_543_47# 0.01fF
C5166 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__dfrtn_1_7/a_193_47# 0.00fF
C5167 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# sky130_fd_sc_hd__dfrtn_1_7/a_27_47# 0.01fF
C5168 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# 0.01fF
C5169 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C5170 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_3/a_448_47# 0.00fF
C5171 DOUT[4] sky130_fd_sc_hd__dfrtn_1_12/a_27_47# 0.00fF
C5172 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__inv_1_0/Y 0.32fF
C5173 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_0/a_651_413# 0.00fF
C5174 sky130_fd_sc_hd__mux4_2_0/a_872_316# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C5175 sky130_fd_sc_hd__dfrtn_1_28/a_193_47# sky130_fd_sc_hd__dfrtn_1_28/a_651_413# -0.00fF
C5176 sky130_fd_sc_hd__dfrtp_1_0/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5177 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C5178 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# VDD 0.01fF
C5179 sky130_fd_sc_hd__dfrtn_1_36/a_761_289# sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C5180 sky130_fd_sc_hd__inv_1_2/A DOUT[8] 0.00fF
C5181 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_31/a_448_47# 0.00fF
C5182 VDD sky130_fd_sc_hd__inv_1_50/Y 0.67fF
C5183 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# 0.00fF
C5184 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__dfrtn_1_6/a_639_47# -0.00fF
C5185 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# DOUT[20] 0.01fF
C5186 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# DOUT[6] 0.00fF
C5187 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C5188 sky130_fd_sc_hd__dfrtn_1_22/a_1108_47# RESET_COUNTERn 0.01fF
C5189 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C5190 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C5191 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_639_47# 0.00fF
C5192 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C5193 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.00fF
C5194 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.01fF
C5195 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# 0.00fF
C5196 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C5197 sky130_fd_sc_hd__dfrtn_1_39/a_651_413# VDD 0.02fF
C5198 sky130_fd_sc_hd__nor3_1_11/a_193_297# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C5199 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_32/a_27_47# 0.02fF
C5200 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5201 CLK_REF sky130_fd_sc_hd__dfrtn_1_20/a_761_289# 0.00fF
C5202 sky130_fd_sc_hd__dfrtn_1_30/a_761_289# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C5203 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_3/a_193_47# 0.00fF
C5204 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_10/a_543_47# -0.00fF
C5205 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_10/a_761_289# -0.00fF
C5206 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__dfrtn_1_3/a_448_47# 0.00fF
C5207 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__dfrtn_1_3/a_1270_413# 0.00fF
C5208 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# sky130_fd_sc_hd__dfrtn_1_3/a_761_289# 0.00fF
C5209 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__dfrtn_1_3/a_543_47# 0.00fF
C5210 sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# sky130_fd_sc_hd__dfrtn_1_3/a_193_47# 0.00fF
C5211 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C5212 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C5213 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C5214 sky130_fd_sc_hd__dfrtn_1_18/a_651_413# VDD 0.01fF
C5215 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C5216 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__dfrtn_1_25/a_448_47# 0.00fF
C5217 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C5218 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C5219 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C5220 sky130_fd_sc_hd__dfrtn_1_41/a_639_47# DOUT[2] 0.00fF
C5221 sky130_fd_sc_hd__dfrtn_1_40/a_1462_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C5222 sky130_fd_sc_hd__dfrtn_1_17/a_543_47# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C5223 sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.01fF
C5224 sky130_fd_sc_hd__dfrtn_1_24/a_1462_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C5225 sky130_fd_sc_hd__dfrtn_1_16/a_543_47# RESET_COUNTERn 0.01fF
C5226 sky130_fd_sc_hd__dfrtn_1_8/a_1283_21# DOUT[21] 0.00fF
C5227 HEADER_2/a_508_138# HEADER_0/a_508_138# 0.00fF
C5228 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# DOUT[14] 0.00fF
C5229 VDD sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.08fF
C5230 sky130_fd_sc_hd__dfrtn_1_9/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5231 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# -0.00fF
C5232 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_20/a_543_47# -0.00fF
C5233 sky130_fd_sc_hd__or3_1_0/X SEL_CONV_TIME[1] 0.14fF
C5234 sky130_fd_sc_hd__nor3_1_19/Y sky130_fd_sc_hd__inv_1_48/A 0.02fF
C5235 outb sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C5236 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C5237 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_639_47# 0.00fF
C5238 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__dfrtn_1_4/a_543_47# 0.00fF
C5239 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C5240 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__nand2_1_1/Y 0.01fF
C5241 sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C5242 sky130_fd_sc_hd__dfrtn_1_41/a_805_47# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C5243 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_805_47# 0.00fF
C5244 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# sky130_fd_sc_hd__dfrtn_1_38/a_639_47# 0.00fF
C5245 sky130_fd_sc_hd__dfrtn_1_19/a_543_47# VDD 0.06fF
C5246 sky130_fd_sc_hd__dfrtp_1_3/a_448_47# DOUT[23] 0.00fF
C5247 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# 0.00fF
C5248 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__dfrtn_1_1/a_27_47# 0.00fF
C5249 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_1/a_543_47# 0.00fF
C5250 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_1/a_639_47# 0.00fF
C5251 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_1/a_448_47# 0.00fF
C5252 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C5253 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# 0.00fF
C5254 sky130_fd_sc_hd__o221ai_1_0/a_109_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5255 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_18/a_543_47# 0.01fF
C5256 sky130_fd_sc_hd__mux4_2_0/a_1060_369# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C5257 sky130_fd_sc_hd__dfrtn_1_24/a_1270_413# SEL_CONV_TIME[1] 0.00fF
C5258 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C5259 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C5260 sky130_fd_sc_hd__dfrtp_1_3/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5261 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_639_47# -0.00fF
C5262 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_33/A 0.21fF
C5263 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.07fF
C5264 sky130_fd_sc_hd__dfrtn_1_16/a_1217_47# DOUT[15] 0.00fF
C5265 sky130_fd_sc_hd__nor3_1_0/a_193_297# DOUT[5] 0.00fF
C5266 sky130_fd_sc_hd__dfrtn_1_33/a_805_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C5267 DOUT[4] sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C5268 sky130_fd_sc_hd__nor3_1_5/a_193_297# DOUT[11] 0.00fF
C5269 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C5270 sky130_fd_sc_hd__dfrtp_1_2/a_448_47# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C5271 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C5272 sky130_fd_sc_hd__dfrtn_1_23/a_1217_47# DOUT[21] 0.00fF
C5273 sky130_fd_sc_hd__dfrtn_1_23/a_448_47# RESET_COUNTERn 0.01fF
C5274 sky130_fd_sc_hd__dfrtn_1_22/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5275 sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C5276 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__or3b_2_0/a_388_297# 0.00fF
C5277 sky130_fd_sc_hd__nor3_1_1/a_109_297# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C5278 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__dfrtn_1_26/a_639_47# 0.00fF
C5279 sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.00fF
C5280 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C5281 sky130_fd_sc_hd__dfrtn_1_12/a_1217_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C5282 sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# DOUT[6] 0.00fF
C5283 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# RESET_COUNTERn 0.01fF
C5284 sky130_fd_sc_hd__dfrtn_1_7/a_448_47# DOUT[20] 0.00fF
C5285 sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# DOUT[7] 0.00fF
C5286 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C5287 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C5288 sky130_fd_sc_hd__inv_1_19/A VIN 0.20fF
C5289 sky130_fd_sc_hd__inv_1_17/A DOUT[10] 0.00fF
C5290 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# -0.00fF
C5291 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# -0.00fF
C5292 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# DOUT[20] 0.00fF
C5293 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# DOUT[7] 0.00fF
C5294 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# RESET_COUNTERn 0.00fF
C5295 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# DOUT[6] 0.00fF
C5296 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# CLK_REF 0.47fF
C5297 DOUT[20] DOUT[8] 0.03fF
C5298 DOUT[6] DOUT[7] 5.14fF
C5299 DOUT[21] RESET_COUNTERn 0.80fF
C5300 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C5301 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__mux4_1_0/a_750_97# -0.00fF
C5302 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_32/a_1217_47# 0.00fF
C5303 sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C5304 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_448_47# 0.00fF
C5305 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# sky130_fd_sc_hd__dfrtn_1_27/a_761_289# 0.00fF
C5306 sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.00fF
C5307 sky130_fd_sc_hd__inv_1_39/A sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C5308 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5309 sky130_fd_sc_hd__o2111a_2_0/a_386_47# sky130_fd_sc_hd__o311a_1_0/a_266_47# 0.00fF
C5310 sky130_fd_sc_hd__dfrtn_1_24/a_651_413# VDD 0.01fF
C5311 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C5312 CLK_REF sky130_fd_sc_hd__dfrtn_1_21/a_639_47# 0.00fF
C5313 sky130_fd_sc_hd__dfrtn_1_16/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5314 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5315 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# VDD 0.04fF
C5316 sky130_fd_sc_hd__dfrtn_1_11/a_805_47# outb 0.00fF
C5317 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5318 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# SEL_CONV_TIME[0] 0.00fF
C5319 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C5320 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_31/a_761_289# 0.00fF
C5321 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__nor3_2_3/B 0.04fF
C5322 sky130_fd_sc_hd__dfrtn_1_9/a_448_47# DOUT[14] 0.00fF
C5323 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__nor3_1_16/a_109_297# 0.00fF
C5324 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C5325 sky130_fd_sc_hd__inv_1_53/A SEL_CONV_TIME[1] 0.08fF
C5326 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C5327 sky130_fd_sc_hd__dfrtn_1_17/a_1462_47# sky130_fd_sc_hd__dfrtn_1_19/a_543_47# 0.00fF
C5328 sky130_fd_sc_hd__dfrtn_1_33/a_761_289# SEL_CONV_TIME[1] 0.00fF
C5329 sky130_fd_sc_hd__dfrtn_1_26/a_805_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C5330 sky130_fd_sc_hd__dfrtn_1_8/a_805_47# RESET_COUNTERn 0.00fF
C5331 sky130_fd_sc_hd__inv_1_1/Y DOUT[9] 0.00fF
C5332 sky130_fd_sc_hd__o311a_1_0/A3 RESET_COUNTERn 0.57fF
C5333 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__or3b_2_0/X 0.01fF
C5334 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# sky130_fd_sc_hd__o211a_1_0/X 0.00fF
C5335 sky130_fd_sc_hd__dfrtn_1_30/a_651_413# SEL_CONV_TIME[1] 0.00fF
C5336 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# DOUT[0] 0.00fF
C5337 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__nor3_1_4/a_193_297# 0.00fF
C5338 sky130_fd_sc_hd__inv_1_28/A sky130_fd_sc_hd__inv_1_28/Y 0.01fF
C5339 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_21/a_27_47# 0.01fF
C5340 sky130_fd_sc_hd__dfrtn_1_32/a_639_47# sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C5341 DOUT[4] sky130_fd_sc_hd__or3b_2_0/a_388_297# 0.00fF
C5342 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5343 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# 0.00fF
C5344 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# 0.00fF
C5345 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# 0.01fF
C5346 sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C5347 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C5348 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C5349 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5350 sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C5351 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C5352 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# VDD 0.04fF
C5353 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C5354 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# sky130_fd_sc_hd__dfrtn_1_23/a_27_47# 0.00fF
C5355 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# SEL_CONV_TIME[1] 0.00fF
C5356 DOUT[4] sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# 0.00fF
C5357 sky130_fd_sc_hd__inv_1_36/A sky130_fd_sc_hd__inv_1_40/A 0.01fF
C5358 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5359 sky130_fd_sc_hd__dfrtn_1_34/a_639_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C5360 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__inv_1_47/Y 0.00fF
C5361 sky130_fd_sc_hd__nor3_2_0/a_281_297# RESET_COUNTERn 0.00fF
C5362 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__dfrtn_1_1/a_448_47# 0.00fF
C5363 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# VDD 0.08fF
C5364 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C5365 sky130_fd_sc_hd__o311a_1_0/a_368_297# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C5366 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__inv_1_40/Y 0.01fF
C5367 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# 0.00fF
C5368 sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5369 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C5370 sky130_fd_sc_hd__dfrtn_1_30/a_448_47# VDD 0.01fF
C5371 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# DOUT[3] 0.01fF
C5372 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__a221oi_4_0/a_453_47# 0.00fF
C5373 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__nor3_1_4/a_109_297# 0.00fF
C5374 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__inv_1_35/A 0.59fF
C5375 sky130_fd_sc_hd__dfrtn_1_16/a_448_47# DOUT[23] 0.00fF
C5376 DOUT[4] sky130_fd_sc_hd__dfrtn_1_31/a_761_289# 0.00fF
C5377 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__inv_1_41/Y 0.02fF
C5378 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C5379 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# DOUT[14] 0.00fF
C5380 sky130_fd_sc_hd__dfrtn_1_14/a_651_413# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C5381 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C5382 sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# CLK_REF 0.00fF
C5383 sky130_fd_sc_hd__inv_1_42/Y SEL_CONV_TIME[1] 0.11fF
C5384 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__dfrtn_1_17/a_543_47# 0.00fF
C5385 sky130_fd_sc_hd__dfrtn_1_14/a_805_47# DOUT[17] 0.00fF
C5386 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_0/a_834_97# -0.00fF
C5387 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_668_97# -0.00fF
C5388 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C5389 sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# sky130_fd_sc_hd__dfrtn_1_27/a_448_47# 0.00fF
C5390 sky130_fd_sc_hd__dfrtn_1_34/a_543_47# SEL_CONV_TIME[1] 0.00fF
C5391 sky130_fd_sc_hd__o211a_1_1/a_215_47# sky130_fd_sc_hd__dfrtn_1_17/a_761_289# 0.00fF
C5392 sky130_fd_sc_hd__o211a_1_1/a_297_297# sky130_fd_sc_hd__dfrtn_1_17/a_543_47# 0.00fF
C5393 sky130_fd_sc_hd__o211a_1_1/a_510_47# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C5394 sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# DOUT[2] 0.00fF
C5395 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C5396 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C5397 sky130_fd_sc_hd__inv_1_42/A sky130_fd_sc_hd__inv_1_48/Y 0.02fF
C5398 sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__o211a_1_0/a_297_297# 0.00fF
C5399 sky130_fd_sc_hd__dfrtn_1_16/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5400 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5401 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__or3b_2_0/B 0.00fF
C5402 sky130_fd_sc_hd__dfrtn_1_8/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5403 sky130_fd_sc_hd__o211a_1_0/a_79_21# sky130_fd_sc_hd__o211a_1_0/a_510_47# -0.00fF
C5404 sky130_fd_sc_hd__dfrtn_1_36/a_1270_413# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C5405 sky130_fd_sc_hd__dfrtn_1_17/a_448_47# sky130_fd_sc_hd__o211a_1_1/X 0.00fF
C5406 sky130_fd_sc_hd__or3_1_0/a_183_297# sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C5407 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C5408 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C5409 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# 0.01fF
C5410 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# sky130_fd_sc_hd__dfrtn_1_11/a_543_47# 0.00fF
C5411 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# 0.00fF
C5412 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__dfrtn_1_11/a_761_289# 0.00fF
C5413 sky130_fd_sc_hd__o211a_1_1/a_297_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5414 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C5415 sky130_fd_sc_hd__o211a_1_1/a_510_47# VDD 0.00fF
C5416 SEL_CONV_TIME[3] DOUT[21] 0.00fF
C5417 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C5418 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# 0.01fF
C5419 VDD sky130_fd_sc_hd__inv_1_36/A 1.26fF
C5420 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_12/a_639_47# 0.00fF
C5421 DOUT[4] sky130_fd_sc_hd__dfrtn_1_32/a_651_413# 0.00fF
C5422 sky130_fd_sc_hd__o2111a_2_0/a_458_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C5423 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_1/a_761_289# -0.00fF
C5424 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C5425 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# sky130_fd_sc_hd__inv_1_6/A 0.23fF
C5426 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__o2111a_2_0/X 0.05fF
C5427 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# 0.00fF
C5428 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# 0.00fF
C5429 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# 0.00fF
C5430 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__dfrtn_1_17/a_651_413# 0.00fF
C5431 sky130_fd_sc_hd__dfrtp_1_2/a_639_47# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C5432 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__dfrtn_1_17/a_543_47# 0.00fF
C5433 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_639_47# 0.00fF
C5434 sky130_fd_sc_hd__dfrtp_1_2/a_805_47# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C5435 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_805_47# 0.00fF
C5436 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__inv_1_8/A 0.01fF
C5437 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# sky130_fd_sc_hd__mux4_1_0/X 0.01fF
C5438 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_14/a_805_47# 0.00fF
C5439 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C5440 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_37/a_193_47# -0.15fF
C5441 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# 0.00fF
C5442 sky130_fd_sc_hd__dfrtp_1_1/D RESET_COUNTERn 0.01fF
C5443 sky130_fd_sc_hd__dfrtn_1_28/a_761_289# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C5444 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__dfrtn_1_42/a_651_413# 0.00fF
C5445 sky130_fd_sc_hd__nor3_2_2/a_281_297# sky130_fd_sc_hd__dfrtn_1_42/a_448_47# 0.00fF
C5446 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# VDD 0.08fF
C5447 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__nor3_2_3/C 0.25fF
C5448 sky130_fd_sc_hd__o211a_1_0/a_297_297# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C5449 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C5450 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# DOUT[14] 0.01fF
C5451 sky130_fd_sc_hd__nor3_1_12/a_193_297# outb 0.00fF
C5452 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5453 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# VDD 0.06fF
C5454 VDD sky130_fd_sc_hd__inv_1_41/Y 0.54fF
C5455 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5456 sky130_fd_sc_hd__dfrtp_1_2/a_639_47# VDD 0.00fF
C5457 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__dfrtn_1_30/a_761_289# 0.00fF
C5458 sky130_fd_sc_hd__or2b_1_0/a_301_297# sky130_fd_sc_hd__dfrtn_1_30/a_27_47# 0.00fF
C5459 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__dfrtn_1_30/a_193_47# 0.00fF
C5460 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_18/a_1217_47# 0.00fF
C5461 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# sky130_fd_sc_hd__inv_1_40/Y 0.13fF
C5462 sky130_fd_sc_hd__dfrtn_1_7/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5463 sky130_fd_sc_hd__dfrtn_1_28/a_761_289# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C5464 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C5465 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C5466 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__inv_1_5/A 0.05fF
C5467 sky130_fd_sc_hd__dfrtn_1_16/a_1108_47# sky130_fd_sc_hd__inv_1_26/A 0.00fF
C5468 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5469 sky130_fd_sc_hd__o311a_1_0/A3 SEL_CONV_TIME[3] 0.01fF
C5470 sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# DOUT[21] 0.01fF
C5471 sky130_fd_sc_hd__dfrtn_1_42/a_1217_47# sky130_fd_sc_hd__dfrtn_1_23/a_27_47# 0.00fF
C5472 sky130_fd_sc_hd__dfrtn_1_12/a_639_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C5473 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C5474 sky130_fd_sc_hd__dfrtn_1_37/a_639_47# RESET_COUNTERn 0.00fF
C5475 sky130_fd_sc_hd__nor3_1_1/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5476 sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# sky130_fd_sc_hd__inv_1_36/A 0.01fF
C5477 sky130_fd_sc_hd__mux4_2_0/a_872_316# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C5478 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C5479 sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# DOUT[3] 0.00fF
C5480 sky130_fd_sc_hd__inv_1_22/A DOUT[12] 0.00fF
C5481 sky130_fd_sc_hd__dfrtn_1_33/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5482 sky130_fd_sc_hd__nor3_1_4/a_109_297# VIN 0.00fF
C5483 sky130_fd_sc_hd__dfrtn_1_33/a_1462_47# VDD -0.00fF
C5484 sky130_fd_sc_hd__dfrtn_1_3/a_1270_413# RESET_COUNTERn 0.00fF
C5485 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__inv_1_43/A 0.07fF
C5486 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C5487 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# HEADER_0/a_508_138# 0.00fF
C5488 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5489 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# VDD 0.07fF
C5490 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# RESET_COUNTERn 0.03fF
C5491 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C5492 sky130_fd_sc_hd__inv_1_54/A SEL_CONV_TIME[0] 0.01fF
C5493 sky130_fd_sc_hd__dfrtn_1_11/a_1270_413# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C5494 SEL_CONV_TIME[2] sky130_fd_sc_hd__o311a_1_0/A3 0.10fF
C5495 SEL_CONV_TIME[0] sky130_fd_sc_hd__inv_1_48/A 0.03fF
C5496 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_10/a_27_47# 0.11fF
C5497 sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# sky130_fd_sc_hd__inv_1_15/A 0.02fF
C5498 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C5499 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C5500 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C5501 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# HEADER_0/a_508_138# 0.00fF
C5502 sky130_fd_sc_hd__dfrtp_1_1/a_448_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C5503 sky130_fd_sc_hd__dfrtn_1_0/a_651_413# DOUT[17] 0.00fF
C5504 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# RESET_COUNTERn 0.16fF
C5505 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# sky130_fd_sc_hd__dfrtn_1_29/a_543_47# 0.00fF
C5506 sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C5507 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# sky130_fd_sc_hd__dfrtn_1_29/a_639_47# 0.00fF
C5508 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# 0.00fF
C5509 sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# sky130_fd_sc_hd__inv_1_28/A 0.01fF
C5510 sky130_fd_sc_hd__nor3_1_3/a_193_297# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C5511 sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# RESET_COUNTERn 0.01fF
C5512 sky130_fd_sc_hd__dfrtn_1_38/a_805_47# VDD 0.00fF
C5513 sky130_fd_sc_hd__dfrtn_1_38/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5514 VDD sky130_fd_sc_hd__inv_1_49/A 0.93fF
C5515 sky130_fd_sc_hd__dfrtn_1_21/a_651_413# RESET_COUNTERn 0.00fF
C5516 sky130_fd_sc_hd__nor3_1_20/a_193_297# DOUT[1] 0.00fF
C5517 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__dfrtn_1_11/a_805_47# 0.00fF
C5518 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C5519 sky130_fd_sc_hd__dfrtn_1_42/a_1270_413# DOUT[15] 0.00fF
C5520 sky130_fd_sc_hd__dfrtn_1_7/a_1462_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C5521 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_40/a_193_47# 0.00fF
C5522 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C5523 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C5524 sky130_fd_sc_hd__dfrtn_1_14/a_761_289# VDD 0.04fF
C5525 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# 0.00fF
C5526 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# sky130_fd_sc_hd__dfrtn_1_0/a_761_289# 0.00fF
C5527 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__dfrtn_1_0/a_543_47# 0.01fF
C5528 sky130_fd_sc_hd__dfrtn_1_12/a_761_289# sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# 0.00fF
C5529 sky130_fd_sc_hd__dfrtn_1_26/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5530 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5531 sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# VDD -0.00fF
C5532 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_0/a_193_47# 0.00fF
C5533 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# DOUT[3] 0.00fF
C5534 sky130_fd_sc_hd__dfrtp_1_0/a_761_289# RESET_COUNTERn 0.01fF
C5535 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_8/Y 0.01fF
C5536 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C5537 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# -0.00fF
C5538 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_41/a_448_47# -0.00fF
C5539 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C5540 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__nor3_1_19/Y 0.05fF
C5541 sky130_fd_sc_hd__dfrtn_1_34/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5542 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5543 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# 0.00fF
C5544 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_8/a_651_413# 0.00fF
C5545 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# lc_out 0.01fF
C5546 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C5547 sky130_fd_sc_hd__dfrtn_1_23/a_1462_47# sky130_fd_sc_hd__inv_1_40/Y 0.00fF
C5548 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_805_47# -0.00fF
C5549 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__inv_1_34/Y 0.01fF
C5550 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C5551 sky130_fd_sc_hd__dfrtn_1_39/a_543_47# RESET_COUNTERn 0.00fF
C5552 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__inv_1_51/Y 0.02fF
C5553 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# sky130_fd_sc_hd__inv_1_39/Y 0.54fF
C5554 sky130_fd_sc_hd__dfrtn_1_25/a_805_47# RESET_COUNTERn 0.00fF
C5555 sky130_fd_sc_hd__nor3_1_11/a_109_297# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C5556 sky130_fd_sc_hd__dfrtp_1_3/a_448_47# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C5557 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# sky130_fd_sc_hd__inv_1_32/Y 0.00fF
C5558 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C5559 sky130_fd_sc_hd__dfrtn_1_18/a_543_47# RESET_COUNTERn 0.00fF
C5560 DOUT[9] RESET_COUNTERn 0.01fF
C5561 sky130_fd_sc_hd__inv_1_42/A sky130_fd_sc_hd__nor3_2_3/B 0.08fF
C5562 sky130_fd_sc_hd__conb_1_0/LO VDD 0.14fF
C5563 sky130_fd_sc_hd__dfrtp_1_0/a_805_47# DOUT[15] 0.00fF
C5564 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# 0.00fF
C5565 DOUT[4] sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# 0.00fF
C5566 sky130_fd_sc_hd__nor3_1_10/a_109_297# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C5567 sky130_fd_sc_hd__dfrtn_1_4/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5568 sky130_fd_sc_hd__or3_1_0/a_183_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5569 en DOUT[6] 0.08fF
C5570 sky130_fd_sc_hd__dfrtn_1_3/a_761_289# sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C5571 sky130_fd_sc_hd__dfrtn_1_28/a_651_413# SEL_CONV_TIME[1] 0.00fF
C5572 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C5573 sky130_fd_sc_hd__dfrtn_1_42/a_1217_47# RESET_COUNTERn 0.00fF
C5574 sky130_fd_sc_hd__mux4_2_0/a_1064_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C5575 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C5576 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# DOUT[3] 0.01fF
C5577 sky130_fd_sc_hd__mux4_2_0/a_1060_369# sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.00fF
C5578 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__o311a_1_0/a_585_47# 0.00fF
C5579 sky130_fd_sc_hd__inv_1_3/Y DOUT[8] 0.01fF
C5580 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# RESET_COUNTERn 0.03fF
C5581 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_10/a_1217_47# 0.00fF
C5582 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C5583 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__mux4_2_0/a_1279_413# -0.00fF
C5584 sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C5585 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# RESET_COUNTERn 0.00fF
C5586 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C5587 CLK_REF sky130_fd_sc_hd__dfrtn_1_17/a_543_47# 0.00fF
C5588 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__inv_1_2/A 0.01fF
C5589 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__inv_1_32/A 0.01fF
C5590 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# SEL_CONV_TIME[0] 0.00fF
C5591 sky130_fd_sc_hd__o221ai_1_0/a_295_297# RESET_COUNTERn 0.00fF
C5592 sky130_fd_sc_hd__nor3_1_17/a_109_297# DOUT[21] 0.00fF
C5593 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__inv_1_36/A 0.01fF
C5594 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__inv_1_42/A 0.02fF
C5595 sky130_fd_sc_hd__inv_1_47/A SEL_CONV_TIME[1] 0.01fF
C5596 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__o2111a_2_0/a_674_297# 0.00fF
C5597 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__dfrtn_1_34/a_639_47# 0.00fF
C5598 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C5599 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__nor3_1_3/a_193_297# 0.00fF
C5600 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_761_289# -0.00fF
C5601 CLK_REF sky130_fd_sc_hd__nor3_2_3/C 0.04fF
C5602 sky130_fd_sc_hd__dfrtn_1_31/a_805_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C5603 sky130_fd_sc_hd__dfrtn_1_35/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_761_289# 0.00fF
C5604 sky130_fd_sc_hd__dfrtn_1_35/a_543_47# sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C5605 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_543_47# 0.00fF
C5606 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_25/a_543_47# -0.00fF
C5607 DOUT[13] sky130_fd_sc_hd__dfrtn_1_31/a_1270_413# 0.00fF
C5608 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# sky130_fd_sc_hd__dfrtn_1_39/a_27_47# 0.00fF
C5609 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# 0.01fF
C5610 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# 0.00fF
C5611 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C5612 sky130_fd_sc_hd__dfrtn_1_37/a_639_47# SEL_CONV_TIME[2] 0.00fF
C5613 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# 0.00fF
C5614 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_7/Y 0.01fF
C5615 sky130_fd_sc_hd__dfrtn_1_28/a_448_47# VDD 0.01fF
C5616 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C5617 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_651_413# -0.00fF
C5618 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_11/a_448_47# -0.00fF
C5619 sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C5620 sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5621 sky130_fd_sc_hd__dfrtn_1_25/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5622 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_37/a_193_47# 0.20fF
C5623 sky130_fd_sc_hd__dfrtn_1_9/a_761_289# sky130_fd_sc_hd__inv_1_12/A 0.03fF
C5624 sky130_fd_sc_hd__inv_1_37/A sky130_fd_sc_hd__nor3_1_4/A 0.03fF
C5625 sky130_fd_sc_hd__or3_1_0/X DOUT[21] 0.01fF
C5626 sky130_fd_sc_hd__dfrtn_1_16/a_543_47# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C5627 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_0/a_1462_47# 0.00fF
C5628 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__dfrtn_1_29/a_651_413# 0.00fF
C5629 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C5630 sky130_fd_sc_hd__dfrtn_1_11/a_761_289# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C5631 sky130_fd_sc_hd__mux4_1_0/a_750_97# SEL_CONV_TIME[1] 0.03fF
C5632 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C5633 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_38/a_543_47# 0.01fF
C5634 sky130_fd_sc_hd__nor3_1_20/a_109_297# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C5635 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C5636 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_6/A 0.44fF
C5637 VDD sky130_fd_sc_hd__inv_1_7/A 2.26fF
C5638 sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C5639 HEADER_1/a_508_138# VIN 0.03fF
C5640 sky130_fd_sc_hd__dfrtn_1_4/a_543_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C5641 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__inv_1_32/Y 0.01fF
C5642 sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# VDD 0.12fF
C5643 sky130_fd_sc_hd__dfrtn_1_22/a_1462_47# sky130_fd_sc_hd__inv_1_39/Y 0.00fF
C5644 sky130_fd_sc_hd__inv_1_18/Y outb 0.01fF
C5645 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C5646 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# RESET_COUNTERn 0.01fF
C5647 sky130_fd_sc_hd__dfrtn_1_24/a_1270_413# DOUT[21] 0.00fF
C5648 sky130_fd_sc_hd__dfrtn_1_42/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5649 sky130_fd_sc_hd__dfrtn_1_25/a_448_47# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C5650 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# DOUT[7] 0.00fF
C5651 CLK_REF sky130_fd_sc_hd__nor3_2_1/a_281_297# 0.00fF
C5652 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__o2111a_2_0/a_566_47# 0.00fF
C5653 DOUT[1] sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.01fF
C5654 sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C5655 sky130_fd_sc_hd__dfrtn_1_20/a_651_413# sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# 0.00fF
C5656 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C5657 sky130_fd_sc_hd__or3_1_0/X sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C5658 sky130_fd_sc_hd__inv_1_26/A DOUT[23] 0.00fF
C5659 sky130_fd_sc_hd__dfrtn_1_23/a_448_47# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C5660 DOUT[1] sky130_fd_sc_hd__inv_1_9/A 0.01fF
C5661 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5662 sky130_fd_sc_hd__dfrtn_1_22/a_448_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C5663 sky130_fd_sc_hd__dfrtn_1_16/a_193_47# DOUT[2] 0.01fF
C5664 sky130_fd_sc_hd__dfrtn_1_42/a_193_47# sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# -0.00fF
C5665 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# sky130_fd_sc_hd__dfrtn_1_42/a_1108_47# -0.00fF
C5666 sky130_fd_sc_hd__dfrtn_1_30/a_1270_413# SEL_CONV_TIME[0] 0.00fF
C5667 sky130_fd_sc_hd__dfrtn_1_25/a_805_47# SEL_CONV_TIME[3] 0.00fF
C5668 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__dfrtn_1_7/a_448_47# 0.00fF
C5669 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C5670 sky130_fd_sc_hd__nor3_1_14/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5671 sky130_fd_sc_hd__mux4_1_0/a_757_363# VDD 0.01fF
C5672 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__inv_1_33/A 0.01fF
C5673 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5674 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C5675 sky130_fd_sc_hd__dfrtn_1_10/a_639_47# VDD 0.00fF
C5676 sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# RESET_COUNTERn 0.00fF
C5677 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_19/a_761_289# 0.00fF
C5678 sky130_fd_sc_hd__nor3_2_2/a_27_297# DOUT[2] 0.01fF
C5679 DOUT[9] sky130_fd_sc_hd__inv_1_7/Y 0.05fF
C5680 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# sky130_fd_sc_hd__dfrtn_1_15/a_27_47# 0.00fF
C5681 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C5682 sky130_fd_sc_hd__dfrtn_1_11/a_761_289# sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# 0.00fF
C5683 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# sky130_fd_sc_hd__dfrtn_1_15/a_193_47# 0.00fF
C5684 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_651_413# 0.00fF
C5685 sky130_fd_sc_hd__dfrtp_1_0/a_1108_47# DOUT[23] 0.00fF
C5686 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_20/a_27_47# 0.01fF
C5687 sky130_fd_sc_hd__o2111a_2_0/a_458_47# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C5688 sky130_fd_sc_hd__dfrtn_1_24/a_1270_413# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C5689 sky130_fd_sc_hd__nor3_1_16/a_109_297# sky130_fd_sc_hd__inv_1_38/A 0.00fF
C5690 sky130_fd_sc_hd__nor3_1_3/a_109_297# DOUT[19] 0.00fF
C5691 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C5692 sky130_fd_sc_hd__dfrtn_1_19/a_805_47# RESET_COUNTERn 0.00fF
C5693 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_543_47# -0.00fF
C5694 sky130_fd_sc_hd__dfrtn_1_27/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_761_289# -0.00fF
C5695 sky130_fd_sc_hd__nor3_1_8/a_193_297# DOUT[8] 0.00fF
C5696 sky130_fd_sc_hd__nor3_1_8/a_109_297# RESET_COUNTERn 0.00fF
C5697 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C5698 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_11/a_761_289# 0.00fF
C5699 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__inv_1_37/A 0.01fF
C5700 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# sky130_fd_sc_hd__inv_1_49/A 0.01fF
C5701 sky130_fd_sc_hd__mux4_2_0/a_193_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C5702 sky130_fd_sc_hd__dfrtn_1_38/a_193_47# SEL_CONV_TIME[0] 0.00fF
C5703 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_448_47# -0.00fF
C5704 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_651_413# -0.00fF
C5705 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# DOUT[6] 0.00fF
C5706 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# DOUT[20] 0.00fF
C5707 sky130_fd_sc_hd__dfrtp_1_0/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5708 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_4/a_448_47# 0.00fF
C5709 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__dfrtn_1_4/a_651_413# 0.00fF
C5710 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C5711 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C5712 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__dfrtn_1_4/a_543_47# 0.00fF
C5713 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C5714 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C5715 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C5716 sky130_fd_sc_hd__dfrtn_1_39/a_543_47# SEL_CONV_TIME[2] 0.00fF
C5717 VDD sky130_fd_sc_hd__inv_1_53/Y 0.14fF
C5718 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__inv_1_44/A 0.01fF
C5719 sky130_fd_sc_hd__dfrtn_1_35/a_639_47# sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# 0.00fF
C5720 sky130_fd_sc_hd__dfrtn_1_35/a_543_47# sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# 0.00fF
C5721 sky130_fd_sc_hd__dfrtn_1_35/a_805_47# sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.00fF
C5722 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# sky130_fd_sc_hd__dfrtn_1_39/a_1217_47# 0.00fF
C5723 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__o211a_1_0/X 0.01fF
C5724 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.00fF
C5725 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__inv_1_45/A 0.00fF
C5726 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__inv_1_2/Y 0.06fF
C5727 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C5728 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C5729 DOUT[1] sky130_fd_sc_hd__dfrtn_1_32/a_27_47# 0.02fF
C5730 sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C5731 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C5732 sky130_fd_sc_hd__dfrtn_1_27/a_651_413# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C5733 sky130_fd_sc_hd__dfrtn_1_12/a_639_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C5734 sky130_fd_sc_hd__dfrtn_1_0/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5735 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_37/a_1462_47# 0.00fF
C5736 sky130_fd_sc_hd__dfrtn_1_35/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5737 sky130_fd_sc_hd__dfrtn_1_0/a_805_47# VDD 0.00fF
C5738 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5739 sky130_fd_sc_hd__dfrtn_1_35/a_448_47# VDD 0.01fF
C5740 sky130_fd_sc_hd__o311a_1_0/a_266_297# SEL_CONV_TIME[1] 0.00fF
C5741 sky130_fd_sc_hd__dfrtn_1_30/a_761_289# RESET_COUNTERn 0.00fF
C5742 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C5743 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__inv_1_15/A 0.00fF
C5744 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C5745 sky130_fd_sc_hd__dfrtn_1_26/a_543_47# SEL_CONV_TIME[0] 0.01fF
C5746 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C5747 sky130_fd_sc_hd__dfrtn_1_3/a_805_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C5748 sky130_fd_sc_hd__mux4_2_0/a_288_47# SEL_CONV_TIME[1] -0.00fF
C5749 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# DOUT[19] 0.01fF
C5750 sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# sky130_fd_sc_hd__or3_1_0/C 0.03fF
C5751 sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# SEL_CONV_TIME[0] 0.00fF
C5752 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C5753 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# VDD 0.05fF
C5754 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_14/a_639_47# 0.00fF
C5755 sky130_fd_sc_hd__dfrtn_1_23/a_651_413# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C5756 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# 0.02fF
C5757 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_24/a_448_47# 0.00fF
C5758 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C5759 sky130_fd_sc_hd__dfrtn_1_39/a_1217_47# sky130_fd_sc_hd__inv_1_32/Y 0.00fF
C5760 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# DONE 0.00fF
C5761 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_448_47# -0.00fF
C5762 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_651_413# -0.00fF
C5763 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# VDD 0.21fF
C5764 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# SLC_0/a_438_293# 0.00fF
C5765 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# SLC_0/a_919_243# 0.00fF
C5766 sky130_fd_sc_hd__dfrtp_1_0/a_761_289# SLC_0/a_264_22# 0.00fF
C5767 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# RESET_COUNTERn 0.00fF
C5768 sky130_fd_sc_hd__dfrtp_1_1/a_805_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C5769 sky130_fd_sc_hd__dfrtp_1_0/a_1283_21# sky130_fd_sc_hd__inv_1_26/A 0.01fF
C5770 sky130_fd_sc_hd__inv_1_53/A sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C5771 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_13/A 0.01fF
C5772 sky130_fd_sc_hd__dfrtn_1_9/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5773 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__nand3b_1_0/a_232_47# 0.00fF
C5774 CLK_REF sky130_fd_sc_hd__dfrtp_1_3/a_448_47# 0.01fF
C5775 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__dfrtn_1_24/a_193_47# 0.00fF
C5776 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C5777 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C5778 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# 0.00fF
C5779 sky130_fd_sc_hd__dfrtn_1_8/a_543_47# outb 0.00fF
C5780 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_12/a_639_47# -0.00fF
C5781 sky130_fd_sc_hd__inv_1_34/Y sky130_fd_sc_hd__or2_2_0/A 0.00fF
C5782 sky130_fd_sc_hd__dfrtn_1_16/a_1462_47# DOUT[2] 0.00fF
C5783 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# 0.00fF
C5784 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_639_47# 0.00fF
C5785 sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# VIN 0.08fF
C5786 sky130_fd_sc_hd__o311a_1_0/a_81_21# VDD 0.13fF
C5787 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfrtn_1_38/a_543_47# 0.00fF
C5788 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_12/a_543_47# 0.00fF
C5789 DOUT[9] sky130_fd_sc_hd__dfrtn_1_4/a_639_47# 0.00fF
C5790 VDD sky130_fd_sc_hd__inv_1_6/Y 0.53fF
C5791 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__inv_1_5/Y 0.04fF
C5792 sky130_fd_sc_hd__mux4_2_0/a_193_369# VDD 0.00fF
C5793 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# out 0.01fF
C5794 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# DOUT[0] 0.00fF
C5795 sky130_fd_sc_hd__dfrtn_1_37/a_1462_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C5796 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C5797 sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C5798 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# VIN 0.00fF
C5799 sky130_fd_sc_hd__inv_1_42/Y DOUT[21] 0.00fF
C5800 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# 0.00fF
C5801 sky130_fd_sc_hd__dfrtn_1_34/a_448_47# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C5802 VIN DOUT[6] 0.19fF
C5803 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_20/a_1217_47# 0.00fF
C5804 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__nor3_2_1/a_27_297# 0.00fF
C5805 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__nor3_2_1/a_281_297# 0.00fF
C5806 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C5807 sky130_fd_sc_hd__o2111a_2_0/a_386_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C5808 sky130_fd_sc_hd__o2111a_2_0/a_80_21# SEL_CONV_TIME[0] 0.01fF
C5809 sky130_fd_sc_hd__dfrtn_1_34/a_543_47# DOUT[21] 0.00fF
C5810 sky130_fd_sc_hd__dfrtn_1_35/a_193_47# sky130_fd_sc_hd__inv_1_38/Y 0.14fF
C5811 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# VDD 0.18fF
C5812 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C5813 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# RESET_COUNTERn 0.03fF
C5814 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C5815 sky130_fd_sc_hd__nor3_1_0/a_193_297# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C5816 sky130_fd_sc_hd__inv_1_45/Y VDD 0.22fF
C5817 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5818 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# VDD 0.06fF
C5819 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C5820 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# DOUT[6] 0.00fF
C5821 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# RESET_COUNTERn 0.00fF
C5822 DOUT[13] SEL_CONV_TIME[0] 0.06fF
C5823 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C5824 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__or3b_2_0/X 0.01fF
C5825 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_34/a_27_47# 0.01fF
C5826 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5827 sky130_fd_sc_hd__nand3b_1_0/a_316_47# VDD 0.00fF
C5828 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__inv_1_45/A 0.00fF
C5829 sky130_fd_sc_hd__o311a_1_0/a_368_297# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C5830 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_1217_47# 0.00fF
C5831 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__dfrtn_1_14/a_448_47# 0.00fF
C5832 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# 0.01fF
C5833 sky130_fd_sc_hd__dfrtn_1_33/a_1270_413# RESET_COUNTERn -0.00fF
C5834 sky130_fd_sc_hd__inv_1_39/Y sky130_fd_sc_hd__nor3_2_3/B 0.24fF
C5835 DOUT[1] sky130_fd_sc_hd__dfrtn_1_32/a_1217_47# 0.00fF
C5836 sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# DOUT[19] 0.00fF
C5837 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__mux4_2_0/a_1281_47# 0.00fF
C5838 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__mux4_2_0/a_1064_47# 0.00fF
C5839 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C5840 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5841 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_18/a_448_47# 0.00fF
C5842 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C5843 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C5844 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# 0.00fF
C5845 sky130_fd_sc_hd__dfrtn_1_3/a_651_413# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.00fF
C5846 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# 0.00fF
C5847 sky130_fd_sc_hd__dfrtn_1_34/a_543_47# sky130_fd_sc_hd__o311a_1_0/A3 0.01fF
C5848 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C5849 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# RESET_COUNTERn 0.24fF
C5850 sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5851 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# sky130_fd_sc_hd__inv_1_31/Y -0.00fF
C5852 sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# sky130_fd_sc_hd__inv_1_34/Y 0.01fF
C5853 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C5854 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# sky130_fd_sc_hd__inv_1_47/A 0.01fF
C5855 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C5856 sky130_fd_sc_hd__dfrtn_1_16/a_639_47# sky130_fd_sc_hd__inv_1_25/A 0.00fF
C5857 sky130_fd_sc_hd__dfrtp_1_0/a_1462_47# SLC_0/a_919_243# 0.00fF
C5858 sky130_fd_sc_hd__dfrtn_1_38/a_448_47# RESET_COUNTERn 0.00fF
C5859 sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C5860 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__o211a_1_1/a_215_47# 0.00fF
C5861 sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# DOUT[18] 0.00fF
C5862 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C5863 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C5864 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_43/A 0.13fF
C5865 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# VDD 0.15fF
C5866 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C5867 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C5868 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C5869 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__dfrtn_1_24/a_1462_47# 0.00fF
C5870 sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C5871 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__or2_2_0/B 0.02fF
C5872 sky130_fd_sc_hd__nor3_1_13/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5873 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# VDD 0.08fF
C5874 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5875 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_10/a_639_47# 0.00fF
C5876 sky130_fd_sc_hd__dfrtn_1_39/a_448_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C5877 sky130_fd_sc_hd__dfrtn_1_17/a_761_289# sky130_fd_sc_hd__inv_1_28/Y 0.01fF
C5878 sky130_fd_sc_hd__inv_1_31/Y sky130_fd_sc_hd__inv_1_32/Y 0.01fF
C5879 sky130_fd_sc_hd__nor3_1_4/A DOUT[14] 0.17fF
C5880 VDD sky130_fd_sc_hd__or3_1_0/C 0.90fF
C5881 sky130_fd_sc_hd__inv_1_7/A DOUT[3] 0.27fF
C5882 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C5883 sky130_fd_sc_hd__mux4_2_0/a_1281_47# VDD 0.00fF
C5884 sky130_fd_sc_hd__mux4_2_0/a_397_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5885 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# DOUT[23] 0.00fF
C5886 sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C5887 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# -0.00fF
C5888 sky130_fd_sc_hd__dfrtn_1_11/a_761_289# DOUT[14] 0.00fF
C5889 sky130_fd_sc_hd__nor3_1_6/a_193_297# DOUT[11] 0.00fF
C5890 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__inv_1_48/Y 0.07fF
C5891 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__o311a_1_0/a_266_47# 0.00fF
C5892 sky130_fd_sc_hd__dfrtn_1_18/a_448_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C5893 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# 0.00fF
C5894 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# sky130_fd_sc_hd__nor3_2_2/A 0.53fF
C5895 sky130_fd_sc_hd__nor3_1_20/a_109_297# DOUT[14] 0.00fF
C5896 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_34/a_193_47# 0.00fF
C5897 sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# RESET_COUNTERn 0.00fF
C5898 sky130_fd_sc_hd__dfrtn_1_37/a_639_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C5899 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C5900 sky130_fd_sc_hd__dfrtn_1_33/a_639_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C5901 VDD sky130_fd_sc_hd__or2b_1_0/X 0.74fF
C5902 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_7/A 0.02fF
C5903 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_3/a_651_413# 0.00fF
C5904 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# sky130_fd_sc_hd__dfrtp_1_3/a_543_47# 0.00fF
C5905 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__dfrtp_1_3/a_761_289# 0.00fF
C5906 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C5907 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_448_47# 0.00fF
C5908 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__o211a_1_0/X 0.00fF
C5909 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C5910 sky130_fd_sc_hd__dfrtn_1_34/a_639_47# RESET_COUNTERn 0.00fF
C5911 sky130_fd_sc_hd__dfrtn_1_33/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5912 sky130_fd_sc_hd__dfrtn_1_16/a_651_413# sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C5913 sky130_fd_sc_hd__dfrtn_1_11/a_1217_47# VDD 0.00fF
C5914 sky130_fd_sc_hd__dfrtn_1_11/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5915 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_21/a_1270_413# 0.00fF
C5916 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_21/a_1217_47# 0.00fF
C5917 sky130_fd_sc_hd__dfrtn_1_19/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_543_47# -0.00fF
C5918 sky130_fd_sc_hd__dfrtn_1_36/a_193_47# sky130_fd_sc_hd__inv_1_40/A 0.01fF
C5919 sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5920 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__dfrtn_1_2/a_448_47# 0.00fF
C5921 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_37/a_543_47# 0.01fF
C5922 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__dfrtn_1_37/a_27_47# 0.00fF
C5923 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_37/a_193_47# 0.00fF
C5924 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_37/a_761_289# 0.00fF
C5925 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# DOUT[2] 0.00fF
C5926 sky130_fd_sc_hd__dfrtn_1_3/a_1462_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C5927 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C5928 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C5929 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_34/a_1217_47# 0.00fF
C5930 sky130_fd_sc_hd__o221ai_1_0/a_109_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# -0.00fF
C5931 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_543_47# 0.00fF
C5932 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.01fF
C5933 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C5934 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__dfrtn_1_2/a_761_289# 0.01fF
C5935 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# 0.01fF
C5936 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__nor3_2_0/A 0.01fF
C5937 sky130_fd_sc_hd__inv_1_15/A DOUT[14] 0.00fF
C5938 sky130_fd_sc_hd__nor3_1_10/a_109_297# DOUT[19] 0.00fF
C5939 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_35/a_448_47# 0.00fF
C5940 sky130_fd_sc_hd__dfrtn_1_34/a_651_413# DONE 0.00fF
C5941 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.01fF
C5942 sky130_fd_sc_hd__dfrtn_1_28/a_1270_413# SEL_CONV_TIME[0] 0.00fF
C5943 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__nor3_2_3/B 0.03fF
C5944 sky130_fd_sc_hd__nor3_1_16/a_109_297# DOUT[4] 0.00fF
C5945 sky130_fd_sc_hd__o211a_1_1/a_215_47# DOUT[23] 0.00fF
C5946 sky130_fd_sc_hd__nor3_1_12/a_109_297# DOUT[12] 0.00fF
C5947 sky130_fd_sc_hd__dfrtn_1_27/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5948 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C5949 DOUT[9] sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C5950 sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.03fF
C5951 sky130_fd_sc_hd__dfrtn_1_27/a_639_47# VDD 0.00fF
C5952 sky130_fd_sc_hd__dfrtp_1_3/a_543_47# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C5953 sky130_fd_sc_hd__dfrtp_1_3/a_761_289# sky130_fd_sc_hd__or2_2_0/a_121_297# 0.00fF
C5954 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__inv_1_31/Y 0.01fF
C5955 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_18/a_639_47# 0.00fF
C5956 DOUT[1] sky130_fd_sc_hd__dfrtn_1_22/a_761_289# 0.00fF
C5957 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__dfrtn_1_1/a_651_413# 0.00fF
C5958 sky130_fd_sc_hd__dfrtn_1_40/a_1462_47# RESET_COUNTERn 0.00fF
C5959 sky130_fd_sc_hd__nor3_1_19/Y sky130_fd_sc_hd__inv_1_44/Y 0.01fF
C5960 sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# sky130_fd_sc_hd__inv_1_45/A 0.00fF
C5961 sky130_fd_sc_hd__nor3_2_3/a_27_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C5962 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_639_47# -0.00fF
C5963 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# DOUT[23] 0.00fF
C5964 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# DOUT[14] 0.00fF
C5965 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_193_47# 0.00fF
C5966 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_27_47# 0.00fF
C5967 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C5968 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C5969 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C5970 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C5971 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C5972 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__nor3_1_0/a_109_297# 0.00fF
C5973 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C5974 VDD DOUT[16] 5.09fF
C5975 sky130_fd_sc_hd__dfrtn_1_36/a_193_47# VDD 0.08fF
C5976 sky130_fd_sc_hd__dfrtn_1_26/a_639_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C5977 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_761_289# 0.00fF
C5978 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_193_47# 0.00fF
C5979 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# SEL_CONV_TIME[3] 0.00fF
C5980 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C5981 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C5982 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# VDD -0.00fF
C5983 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C5984 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_5/a_805_47# 0.00fF
C5985 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# 0.00fF
C5986 sky130_fd_sc_hd__dfrtn_1_0/a_543_47# sky130_fd_sc_hd__nor3_1_0/A 0.02fF
C5987 sky130_fd_sc_hd__dfrtn_1_17/a_193_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C5988 sky130_fd_sc_hd__nor3_2_3/C DOUT[12] 0.04fF
C5989 sky130_fd_sc_hd__dfrtp_1_3/a_1217_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C5990 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# 0.00fF
C5991 sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C5992 sky130_fd_sc_hd__dfrtn_1_34/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C5993 sky130_fd_sc_hd__dfrtn_1_12/a_1462_47# VDD 0.00fF
C5994 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_30/a_805_47# 0.00fF
C5995 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_1/a_448_47# 0.00fF
C5996 sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__dfrtn_1_16/a_27_47# 0.00fF
C5997 sky130_fd_sc_hd__dfrtn_1_14/a_448_47# sky130_fd_sc_hd__nor3_1_1/a_109_297# 0.00fF
C5998 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# sky130_fd_sc_hd__nor3_1_1/a_193_297# 0.00fF
C5999 DOUT[4] sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C6000 sky130_fd_sc_hd__dfrtn_1_28/a_651_413# DOUT[21] 0.00fF
C6001 sky130_fd_sc_hd__dfrtn_1_28/a_761_289# RESET_COUNTERn 0.01fF
C6002 sky130_fd_sc_hd__dfrtn_1_33/a_1217_47# DOUT[23] 0.00fF
C6003 sky130_fd_sc_hd__inv_1_38/A sky130_fd_sc_hd__inv_1_36/A 0.00fF
C6004 sky130_fd_sc_hd__dfrtn_1_39/a_543_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C6005 sky130_fd_sc_hd__dfrtn_1_30/a_543_47# sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C6006 VDD sky130_fd_sc_hd__or2_2_0/A 0.36fF
C6007 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# DOUT[9] 0.00fF
C6008 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_21/a_1462_47# 0.00fF
C6009 sky130_fd_sc_hd__dfrtn_1_14/a_639_47# RESET_COUNTERn 0.00fF
C6010 sky130_fd_sc_hd__mux4_1_0/a_1290_413# SEL_CONV_TIME[0] 0.00fF
C6011 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_11/a_27_47# 0.00fF
C6012 sky130_fd_sc_hd__dfrtn_1_42/a_1217_47# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C6013 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_34/a_1462_47# 0.00fF
C6014 DOUT[19] sky130_fd_sc_hd__inv_1_6/A 0.03fF
C6015 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_4/Y 0.24fF
C6016 sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# sky130_fd_sc_hd__dfrtp_1_3/a_651_413# 0.00fF
C6017 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# SEL_CONV_TIME[2] 0.01fF
C6018 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# VIN 0.00fF
C6019 sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C6020 sky130_fd_sc_hd__dfrtn_1_32/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.00fF
C6021 sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C6022 sky130_fd_sc_hd__dfrtn_1_4/a_448_47# VIN 0.00fF
C6023 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C6024 sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# DOUT[22] 0.00fF
C6025 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C6026 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C6027 sky130_fd_sc_hd__inv_1_7/A DOUT[20] 0.04fF
C6028 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C6029 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C6030 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C6031 sky130_fd_sc_hd__inv_1_47/A DOUT[21] 0.00fF
C6032 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__dfrtn_1_37/a_448_47# 0.00fF
C6033 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# 0.00fF
C6034 sky130_fd_sc_hd__dfrtn_1_32/a_193_47# sky130_fd_sc_hd__inv_1_9/A 0.27fF
C6035 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# RESET_COUNTERn 0.03fF
C6036 sky130_fd_sc_hd__inv_1_6/Y DOUT[3] 0.00fF
C6037 sky130_fd_sc_hd__dfrtn_1_18/a_193_47# DOUT[2] 0.03fF
C6038 DOUT[1] sky130_fd_sc_hd__dfrtn_1_23/a_543_47# 0.00fF
C6039 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C6040 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_25/a_448_47# 0.00fF
C6041 sky130_fd_sc_hd__dfrtn_1_22/a_651_413# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C6042 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_24/a_805_47# -0.00fF
C6043 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# -0.00fF
C6044 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_6/Y 0.01fF
C6045 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# -0.23fF
C6046 sky130_fd_sc_hd__o2111a_2_0/a_458_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6047 sky130_fd_sc_hd__dfrtn_1_42/a_639_47# DOUT[2] 0.00fF
C6048 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_3/A 0.03fF
C6049 sky130_fd_sc_hd__o221ai_1_0/a_109_47# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C6050 sky130_fd_sc_hd__nor3_1_12/a_109_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6051 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.03fF
C6052 sky130_fd_sc_hd__or3b_2_0/a_472_297# VDD 0.00fF
C6053 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_448_47# -0.00fF
C6054 sky130_fd_sc_hd__dfrtn_1_31/a_1283_21# SEL_CONV_TIME[1] 0.00fF
C6055 sky130_fd_sc_hd__mux4_1_0/a_193_413# RESET_COUNTERn 0.00fF
C6056 sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# RESET_COUNTERn -0.00fF
C6057 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_41/a_639_47# 0.00fF
C6058 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__o311a_1_0/A3 0.02fF
C6059 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_19/a_448_47# 0.00fF
C6060 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_31/a_761_289# 0.00fF
C6061 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_193_47# 0.00fF
C6062 sky130_fd_sc_hd__or3b_2_0/a_388_297# sky130_fd_sc_hd__dfrtn_1_31/a_27_47# 0.00fF
C6063 sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# DOUT[23] 0.00fF
C6064 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# DOUT[19] 0.00fF
C6065 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# 0.00fF
C6066 sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C6067 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# 0.00fF
C6068 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# 0.00fF
C6069 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C6070 sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# VDD 0.07fF
C6071 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.06fF
C6072 sky130_fd_sc_hd__dfrtn_1_25/a_805_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C6073 sky130_fd_sc_hd__dfrtn_1_17/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6074 SLC_0/a_438_293# outb 0.00fF
C6075 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C6076 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__inv_1_54/Y 0.00fF
C6077 sky130_fd_sc_hd__dfrtn_1_3/a_651_413# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C6078 sky130_fd_sc_hd__dfrtn_1_36/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6079 sky130_fd_sc_hd__dfrtn_1_14/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6080 sky130_fd_sc_hd__dfrtn_1_36/a_1462_47# VDD 0.00fF
C6081 sky130_fd_sc_hd__dfrtn_1_32/a_27_47# sky130_fd_sc_hd__dfrtn_1_32/a_193_47# -0.03fF
C6082 sky130_fd_sc_hd__nor3_1_20/a_109_297# sky130_fd_sc_hd__dfrtn_1_22/a_1283_21# 0.00fF
C6083 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# 0.00fF
C6084 sky130_fd_sc_hd__dfrtn_1_12/a_639_47# sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# 0.00fF
C6085 DOUT[9] sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C6086 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__o2111a_2_0/a_458_47# 0.00fF
C6087 sky130_fd_sc_hd__dfrtn_1_40/a_1462_47# SEL_CONV_TIME[3] 0.00fF
C6088 sky130_fd_sc_hd__nor3_1_4/a_193_297# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C6089 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__o2111a_2_0/a_458_47# 0.00fF
C6090 sky130_fd_sc_hd__nor3_2_3/a_281_297# sky130_fd_sc_hd__dfrtn_1_42/a_448_47# 0.00fF
C6091 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_13/a_651_413# 0.00fF
C6092 sky130_fd_sc_hd__dfrtn_1_17/a_1462_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C6093 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# sky130_fd_sc_hd__inv_1_37/A 0.02fF
C6094 DOUT[1] DOUT[15] 0.00fF
C6095 sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C6096 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C6097 sky130_fd_sc_hd__nor3_1_7/a_109_297# DOUT[14] 0.00fF
C6098 sky130_fd_sc_hd__nor3_2_1/A DOUT[15] 0.58fF
C6099 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.01fF
C6100 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.01fF
C6101 sky130_fd_sc_hd__o311a_1_0/a_585_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C6102 sky130_fd_sc_hd__o211a_1_1/a_510_47# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C6103 sky130_fd_sc_hd__o211a_1_0/a_215_47# DOUT[15] 0.00fF
C6104 sky130_fd_sc_hd__o311a_1_0/a_368_297# SEL_CONV_TIME[0] 0.00fF
C6105 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6106 sky130_fd_sc_hd__dfrtn_1_31/a_543_47# VDD 0.07fF
C6107 sky130_fd_sc_hd__mux4_2_0/a_600_345# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C6108 sky130_fd_sc_hd__mux4_2_0/a_372_413# SEL_CONV_TIME[0] 0.00fF
C6109 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_11/a_1217_47# 0.00fF
C6110 sky130_fd_sc_hd__dfrtn_1_0/a_448_47# RESET_COUNTERn 0.00fF
C6111 sky130_fd_sc_hd__dfrtn_1_35/a_761_289# RESET_COUNTERn 0.02fF
C6112 sky130_fd_sc_hd__dfrtn_1_35/a_651_413# DOUT[21] 0.00fF
C6113 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_1_19/A 0.00fF
C6114 sky130_fd_sc_hd__nor3_1_11/a_109_297# sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# 0.00fF
C6115 sky130_fd_sc_hd__dfrtn_1_3/a_805_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C6116 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__dfrtn_1_28/a_27_47# 0.00fF
C6117 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# sky130_fd_sc_hd__or2b_1_0/X 0.01fF
C6118 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_761_289# -0.00fF
C6119 sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__nor3_2_3/B 0.07fF
C6120 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C6121 sky130_fd_sc_hd__or2b_1_0/a_27_53# SEL_CONV_TIME[1] 0.02fF
C6122 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# DOUT[3] 0.00fF
C6123 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__dfrtn_1_39/a_27_47# 0.00fF
C6124 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_39/a_543_47# 0.00fF
C6125 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_1270_413# 0.00fF
C6126 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_639_47# 0.00fF
C6127 sky130_fd_sc_hd__dfrtn_1_40/a_1462_47# SEL_CONV_TIME[2] 0.00fF
C6128 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_30/a_448_47# 0.00fF
C6129 sky130_fd_sc_hd__nor3_1_4/a_193_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6130 sky130_fd_sc_hd__dfrtn_1_32/a_1462_47# sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.00fF
C6131 sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# sky130_fd_sc_hd__dfrtn_1_36/a_1462_47# 0.00fF
C6132 sky130_fd_sc_hd__inv_1_8/Y RESET_COUNTERn 0.28fF
C6133 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C6134 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C6135 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C6136 sky130_fd_sc_hd__dfrtn_1_32/a_1462_47# sky130_fd_sc_hd__inv_1_9/A 0.00fF
C6137 sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# DOUT[22] 0.00fF
C6138 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__inv_1_31/A 0.00fF
C6139 sky130_fd_sc_hd__dfrtn_1_20/a_1217_47# RESET_COUNTERn -0.00fF
C6140 sky130_fd_sc_hd__dfrtn_1_41/a_651_413# SEL_CONV_TIME[0] 0.00fF
C6141 sky130_fd_sc_hd__inv_1_45/A VDD 0.76fF
C6142 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__inv_1_43/Y 0.02fF
C6143 sky130_fd_sc_hd__or2_2_0/B DOUT[15] 0.01fF
C6144 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# sky130_fd_sc_hd__o221ai_1_0/a_493_297# 0.00fF
C6145 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C6146 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C6147 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.01fF
C6148 sky130_fd_sc_hd__dfrtp_1_2/a_639_47# sky130_fd_sc_hd__inv_1_29/Y 0.00fF
C6149 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_2/A 0.02fF
C6150 sky130_fd_sc_hd__dfrtn_1_18/a_1462_47# DOUT[2] 0.00fF
C6151 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_18/a_543_47# 0.00fF
C6152 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C6153 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_1270_413# 0.00fF
C6154 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_18/a_761_289# 0.00fF
C6155 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_639_47# 0.00fF
C6156 sky130_fd_sc_hd__inv_1_33/Y VDD 0.72fF
C6157 sky130_fd_sc_hd__dfrtn_1_42/a_448_47# sky130_fd_sc_hd__inv_1_25/A 0.00fF
C6158 sky130_fd_sc_hd__dfrtn_1_32/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6159 sky130_fd_sc_hd__dfrtn_1_32/a_1270_413# VDD 0.00fF
C6160 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6161 sky130_fd_sc_hd__dfrtn_1_7/a_543_47# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C6162 sky130_fd_sc_hd__nor3_2_1/a_281_297# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C6163 sky130_fd_sc_hd__dfrtn_1_4/a_448_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C6164 sky130_fd_sc_hd__dfrtn_1_36/a_651_413# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C6165 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_1/a_193_47# -0.07fF
C6166 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_38/a_639_47# 0.00fF
C6167 sky130_fd_sc_hd__dfrtn_1_36/a_448_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C6168 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C6169 sky130_fd_sc_hd__o311a_1_0/a_266_297# DOUT[21] 0.00fF
C6170 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C6171 sky130_fd_sc_hd__dfrtp_1_3/a_1283_21# sky130_fd_sc_hd__or2_2_0/A 0.01fF
C6172 sky130_fd_sc_hd__inv_1_6/Y DOUT[20] 0.01fF
C6173 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# SEL_CONV_TIME[0] 0.00fF
C6174 sky130_fd_sc_hd__or2b_1_0/a_219_297# VDD 0.05fF
C6175 sky130_fd_sc_hd__mux4_1_0/a_834_97# RESET_COUNTERn 0.01fF
C6176 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_26/a_651_413# 0.00fF
C6177 sky130_fd_sc_hd__dfrtn_1_23/a_761_289# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C6178 sky130_fd_sc_hd__o2111a_2_0/a_458_47# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C6179 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_24/a_651_413# 0.00fF
C6180 sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# sky130_fd_sc_hd__dfrtn_1_28/a_193_47# 0.00fF
C6181 sky130_fd_sc_hd__inv_1_10/A DOUT[16] 0.00fF
C6182 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.02fF
C6183 sky130_fd_sc_hd__nor3_1_15/a_109_297# sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C6184 sky130_fd_sc_hd__nor3_1_12/a_193_297# sky130_fd_sc_hd__inv_1_9/Y 0.00fF
C6185 sky130_fd_sc_hd__o211a_1_0/a_510_47# lc_out 0.00fF
C6186 sky130_fd_sc_hd__dfrtn_1_28/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6187 sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C6188 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__inv_1_14/A 0.15fF
C6189 sky130_fd_sc_hd__nand2_1_1/a_113_47# SEL_CONV_TIME[0] 0.00fF
C6190 sky130_fd_sc_hd__dfrtn_1_4/a_761_289# DOUT[11] 0.00fF
C6191 sky130_fd_sc_hd__dfrtn_1_0/a_651_413# sky130_fd_sc_hd__nor3_1_0/a_193_297# 0.00fF
C6192 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C6193 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C6194 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# VDD 0.07fF
C6195 sky130_fd_sc_hd__inv_1_12/A sky130_fd_sc_hd__inv_1_13/A 0.00fF
C6196 sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6197 sky130_fd_sc_hd__dfrtn_1_14/a_543_47# DOUT[9] 0.00fF
C6198 sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C6199 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__inv_1_33/A 0.01fF
C6200 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# RESET_COUNTERn 0.02fF
C6201 sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# 0.00fF
C6202 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_34/a_761_289# 0.00fF
C6203 sky130_fd_sc_hd__dfrtn_1_22/a_1462_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C6204 sky130_fd_sc_hd__o311a_1_0/a_266_297# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C6205 DOUT[4] sky130_fd_sc_hd__dfrtn_1_30/a_448_47# 0.00fF
C6206 sky130_fd_sc_hd__o221ai_1_0/a_493_297# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C6207 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_639_47# 0.00fF
C6208 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C6209 sky130_fd_sc_hd__dfrtn_1_19/a_543_47# sky130_fd_sc_hd__inv_1_28/A 0.02fF
C6210 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfrtn_1_41/a_639_47# 0.00fF
C6211 sky130_fd_sc_hd__nand2_1_0/a_113_47# VIN 0.00fF
C6212 sky130_fd_sc_hd__dfrtn_1_3/a_761_289# sky130_fd_sc_hd__inv_1_8/Y 0.01fF
C6213 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C6214 sky130_fd_sc_hd__dfrtn_1_3/a_639_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C6215 sky130_fd_sc_hd__dfrtn_1_38/a_639_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C6216 sky130_fd_sc_hd__dfrtn_1_28/a_639_47# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C6217 sky130_fd_sc_hd__dfrtn_1_25/a_448_47# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C6218 sky130_fd_sc_hd__dfrtn_1_32/a_761_289# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C6219 sky130_fd_sc_hd__inv_1_34/A DOUT[2] 0.00fF
C6220 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__o211a_1_1/X 0.01fF
C6221 sky130_fd_sc_hd__inv_1_1/Y VDD 0.53fF
C6222 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C6223 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_1/a_761_289# 0.00fF
C6224 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C6225 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# DOUT[3] 0.00fF
C6226 SEL_CONV_TIME[0] sky130_fd_sc_hd__inv_1_44/Y 0.13fF
C6227 sky130_fd_sc_hd__dfrtp_1_1/a_805_47# RESET_COUNTERn 0.00fF
C6228 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__dfrtn_1_25/a_27_47# 0.00fF
C6229 sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__dfrtn_1_25/a_193_47# 0.00fF
C6230 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_25/a_761_289# 0.00fF
C6231 sky130_fd_sc_hd__dfrtp_1_3/a_1108_47# sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# 0.00fF
C6232 sky130_fd_sc_hd__dfrtp_1_3/a_639_47# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C6233 sky130_fd_sc_hd__dfrtp_1_3/a_448_47# sky130_fd_sc_hd__dfrtn_1_17/a_543_47# 0.00fF
C6234 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_639_47# 0.00fF
C6235 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C6236 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# sky130_fd_sc_hd__nor3_1_0/A 0.01fF
C6237 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C6238 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtp_1_2/a_543_47# -0.00fF
C6239 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C6240 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C6241 sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6242 DOUT[4] sky130_fd_sc_hd__inv_1_36/A 0.00fF
C6243 sky130_fd_sc_hd__inv_1_22/A en 0.00fF
C6244 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__inv_1_7/A 0.01fF
C6245 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# 0.00fF
C6246 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__dfrtn_1_29/a_448_47# 0.00fF
C6247 sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# sky130_fd_sc_hd__inv_1_7/A 0.02fF
C6248 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__nor3_1_19/Y 0.03fF
C6249 sky130_fd_sc_hd__o211a_1_0/a_510_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6250 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__dfrtn_1_24/a_193_47# 0.00fF
C6251 sky130_fd_sc_hd__inv_1_34/Y RESET_COUNTERn 0.08fF
C6252 sky130_fd_sc_hd__dfrtp_1_3/a_1270_413# VDD 0.00fF
C6253 sky130_fd_sc_hd__dfrtp_1_3/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6254 DOUT[13] sky130_fd_sc_hd__inv_1_36/Y 0.02fF
C6255 sky130_fd_sc_hd__dfrtn_1_29/a_805_47# SEL_CONV_TIME[1] 0.00fF
C6256 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C6257 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__inv_1_49/A 0.03fF
C6258 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C6259 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__dfrtn_1_24/a_27_47# 0.00fF
C6260 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__dfrtn_1_24/a_193_47# 0.00fF
C6261 sky130_fd_sc_hd__dfrtn_1_28/a_193_47# sky130_fd_sc_hd__inv_1_48/A 0.23fF
C6262 sky130_fd_sc_hd__dfrtn_1_27/a_1217_47# SEL_CONV_TIME[0] 0.00fF
C6263 DOUT[4] sky130_fd_sc_hd__dfrtn_1_34/a_761_289# 0.01fF
C6264 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# sky130_fd_sc_hd__dfrtp_1_1/D 0.00fF
C6265 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__o211a_1_1/a_215_47# 0.00fF
C6266 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_36/a_1462_47# 0.00fF
C6267 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__inv_1_40/A 0.01fF
C6268 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_448_47# -0.00fF
C6269 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# -0.00fF
C6270 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# RESET_COUNTERn 0.01fF
C6271 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_10/a_761_289# 0.01fF
C6272 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# DOUT[23] 0.00fF
C6273 sky130_fd_sc_hd__dfrtn_1_35/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6274 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# DOUT[19] 0.00fF
C6275 sky130_fd_sc_hd__nor3_1_15/a_193_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6276 sky130_fd_sc_hd__dfrtn_1_8/a_761_289# DOUT[12] 0.00fF
C6277 sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# RESET_COUNTERn 0.00fF
C6278 sky130_fd_sc_hd__nor3_1_11/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6279 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C6280 sky130_fd_sc_hd__dfrtn_1_29/a_639_47# VDD 0.00fF
C6281 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__inv_1_53/A 0.02fF
C6282 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# -0.25fF
C6283 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C6284 sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6285 CLK_REF sky130_fd_sc_hd__dfrtn_1_19/a_761_289# 0.01fF
C6286 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__o211a_1_1/a_215_47# 0.00fF
C6287 sky130_fd_sc_hd__dfrtp_1_2/a_639_47# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.00fF
C6288 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C6289 sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# sky130_fd_sc_hd__dfrtn_1_18/a_543_47# 0.00fF
C6290 sky130_fd_sc_hd__dfrtn_1_20/a_1270_413# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C6291 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C6292 sky130_fd_sc_hd__dfrtn_1_18/a_193_47# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C6293 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C6294 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C6295 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_34/a_761_289# 0.00fF
C6296 sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# sky130_fd_sc_hd__inv_1_46/Y 0.01fF
C6297 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__o211a_1_0/a_79_21# 0.01fF
C6298 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__o211a_1_0/a_297_297# 0.00fF
C6299 sky130_fd_sc_hd__dfrtn_1_23/a_651_413# sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C6300 sky130_fd_sc_hd__dfrtn_1_23/a_1270_413# sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C6301 sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# sky130_fd_sc_hd__dfrtn_1_36/a_543_47# 0.00fF
C6302 sky130_fd_sc_hd__dfrtn_1_23/a_761_289# sky130_fd_sc_hd__dfrtn_1_36/a_448_47# 0.00fF
C6303 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C6304 sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# RESET_COUNTERn 0.02fF
C6305 sky130_fd_sc_hd__dfrtn_1_27/a_805_47# DOUT[21] 0.00fF
C6306 sky130_fd_sc_hd__dfrtn_1_38/a_448_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C6307 sky130_fd_sc_hd__dfrtn_1_35/a_448_47# sky130_fd_sc_hd__inv_1_38/A 0.00fF
C6308 sky130_fd_sc_hd__nor3_1_18/a_109_297# RESET_COUNTERn 0.00fF
C6309 sky130_fd_sc_hd__dfrtn_1_11/a_639_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C6310 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C6311 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C6312 DOUT[4] sky130_fd_sc_hd__inv_1_49/A 0.06fF
C6313 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# VDD 0.20fF
C6314 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_25/a_805_47# 0.00fF
C6315 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__dfrtn_1_25/a_639_47# 0.00fF
C6316 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_32/a_1270_413# 0.00fF
C6317 sky130_fd_sc_hd__dfrtn_1_30/a_543_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C6318 sky130_fd_sc_hd__nor3_2_0/a_281_297# sky130_fd_sc_hd__dfrtn_1_12/a_761_289# 0.00fF
C6319 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__dfrtn_1_34/a_193_47# -0.00fF
C6320 DOUT[13] sky130_fd_sc_hd__dfrtn_1_30/a_193_47# 0.02fF
C6321 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C6322 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C6323 sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# DOUT[2] 0.00fF
C6324 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# sky130_fd_sc_hd__mux4_2_0/a_872_316# 0.00fF
C6325 sky130_fd_sc_hd__dfrtn_1_37/a_639_47# sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.00fF
C6326 sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C6327 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# sky130_fd_sc_hd__mux4_2_0/a_193_47# 0.00fF
C6328 sky130_fd_sc_hd__mux4_2_0/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6329 sky130_fd_sc_hd__dfrtn_1_10/a_639_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C6330 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_1283_21# 0.00fF
C6331 sky130_fd_sc_hd__dfrtn_1_36/a_761_289# DOUT[21] 0.00fF
C6332 sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C6333 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# sky130_fd_sc_hd__inv_1_32/A 0.03fF
C6334 sky130_fd_sc_hd__dfrtn_1_21/a_1270_413# VDD 0.00fF
C6335 sky130_fd_sc_hd__nor3_2_3/a_27_297# DOUT[2] 0.00fF
C6336 sky130_fd_sc_hd__o221ai_1_0/a_295_297# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C6337 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# RESET_COUNTERn 0.01fF
C6338 sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C6339 sky130_fd_sc_hd__dfrtn_1_33/a_448_47# sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# 0.00fF
C6340 sky130_fd_sc_hd__dfrtn_1_14/a_761_289# sky130_fd_sc_hd__inv_1_0/Y 0.01fF
C6341 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C6342 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C6343 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__nor3_1_1/a_193_297# 0.00fF
C6344 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# sky130_fd_sc_hd__nor3_1_1/a_109_297# 0.00fF
C6345 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# VDD 0.04fF
C6346 sky130_fd_sc_hd__dfrtn_1_22/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6347 sky130_fd_sc_hd__dfrtn_1_4/a_651_413# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C6348 sky130_fd_sc_hd__dfrtn_1_22/a_805_47# VDD 0.00fF
C6349 DOUT[1] sky130_fd_sc_hd__dfrtn_1_42/a_1270_413# 0.00fF
C6350 sky130_fd_sc_hd__nor3_1_12/a_109_297# sky130_fd_sc_hd__dfrtn_1_8/a_761_289# 0.00fF
C6351 sky130_fd_sc_hd__nor3_1_12/a_193_297# sky130_fd_sc_hd__dfrtn_1_8/a_193_47# 0.00fF
C6352 sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6353 sky130_fd_sc_hd__dfrtn_1_12/a_1270_413# RESET_COUNTERn -0.00fF
C6354 sky130_fd_sc_hd__dfrtn_1_38/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# -0.00fF
C6355 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_448_47# -0.00fF
C6356 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_1/A 0.02fF
C6357 sky130_fd_sc_hd__dfrtn_1_28/a_1462_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C6358 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__dfrtn_1_21/a_193_47# -0.04fF
C6359 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__dfrtn_1_25/a_761_289# 0.00fF
C6360 sky130_fd_sc_hd__nand3b_1_0/a_316_47# sky130_fd_sc_hd__dfrtn_1_25/a_27_47# 0.00fF
C6361 sky130_fd_sc_hd__nand3b_1_0/a_232_47# sky130_fd_sc_hd__dfrtn_1_25/a_193_47# 0.00fF
C6362 sky130_fd_sc_hd__dfrtn_1_26/a_448_47# DOUT[2] 0.00fF
C6363 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# 0.00fF
C6364 sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# 0.00fF
C6365 sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# sky130_fd_sc_hd__dfrtn_1_34/a_1462_47# 0.00fF
C6366 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__inv_1_28/Y 0.04fF
C6367 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# 0.00fF
C6368 sky130_fd_sc_hd__inv_1_37/A sky130_fd_sc_hd__nor3_2_3/B 0.54fF
C6369 sky130_fd_sc_hd__nor3_1_11/a_193_297# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C6370 sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# sky130_fd_sc_hd__inv_1_53/Y 0.01fF
C6371 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__dfrtn_1_6/a_448_47# 0.00fF
C6372 sky130_fd_sc_hd__dfrtn_1_23/a_1217_47# sky130_fd_sc_hd__inv_1_40/A 0.00fF
C6373 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# 0.00fF
C6374 sky130_fd_sc_hd__dfrtp_1_0/a_761_289# sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# 0.00fF
C6375 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# sky130_fd_sc_hd__dfrtp_1_1/a_27_47# 0.00fF
C6376 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# 0.00fF
C6377 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C6378 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__inv_1_49/A 0.00fF
C6379 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# 0.00fF
C6380 sky130_fd_sc_hd__inv_1_52/A DOUT[1] 0.02fF
C6381 sky130_fd_sc_hd__dfrtn_1_0/a_1270_413# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C6382 sky130_fd_sc_hd__dfrtn_1_8/a_1270_413# sky130_fd_sc_hd__inv_1_9/A 0.00fF
C6383 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__nor3_1_4/a_109_297# 0.00fF
C6384 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__nor3_1_4/A 0.01fF
C6385 sky130_fd_sc_hd__dfrtn_1_26/a_543_47# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C6386 sky130_fd_sc_hd__dfrtn_1_27/a_448_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C6387 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_1270_413# 0.00fF
C6388 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C6389 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C6390 sky130_fd_sc_hd__mux4_2_0/a_1060_369# SEL_CONV_TIME[3] 0.00fF
C6391 sky130_fd_sc_hd__dfrtn_1_3/a_805_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C6392 sky130_fd_sc_hd__dfrtn_1_16/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C6393 sky130_fd_sc_hd__dfrtn_1_27/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C6394 sky130_fd_sc_hd__dfrtn_1_16/a_1270_413# VDD 0.00fF
C6395 sky130_fd_sc_hd__dfrtn_1_8/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C6396 sky130_fd_sc_hd__dfrtn_1_8/a_1283_21# VDD 0.11fF
C6397 sky130_fd_sc_hd__nor3_1_3/a_193_297# DOUT[14] 0.00fF
C6398 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_543_47# -0.00fF
C6399 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__dfrtn_1_29/a_761_289# -0.00fF
C6400 sky130_fd_sc_hd__dfrtn_1_40/a_1462_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C6401 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_1217_47# -0.00fF
C6402 sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C6403 sky130_fd_sc_hd__a221oi_4_0/a_27_297# RESET_COUNTERn 0.00fF
C6404 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C6405 sky130_fd_sc_hd__inv_1_40/A RESET_COUNTERn 0.27fF
C6406 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C6407 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_20/a_448_47# 0.00fF
C6408 sky130_fd_sc_hd__nor3_1_13/a_193_297# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C6409 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C6410 sky130_fd_sc_hd__dfrtn_1_31/a_1108_47# SEL_CONV_TIME[0] 0.01fF
C6411 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C6412 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_40/a_448_47# -0.00fF
C6413 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_40/a_651_413# -0.00fF
C6414 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# DOUT[2] 0.00fF
C6415 sky130_fd_sc_hd__dfrtp_1_0/a_805_47# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C6416 sky130_fd_sc_hd__inv_1_3/A DOUT[7] 0.03fF
C6417 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C6418 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C6419 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6420 sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C6421 sky130_fd_sc_hd__mux4_2_0/a_1060_369# SEL_CONV_TIME[2] 0.00fF
C6422 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__or3_1_0/C 0.05fF
C6423 sky130_fd_sc_hd__dfrtn_1_23/a_1217_47# VDD 0.00fF
C6424 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6425 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__conb_1_0/LO 0.00fF
C6426 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__nor3_2_3/B 1.09fF
C6427 DOUT[13] sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# 0.00fF
C6428 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.06fF
C6429 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_1462_47# 0.00fF
C6430 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# 0.00fF
C6431 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C6432 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__or3b_2_0/a_27_47# 0.00fF
C6433 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# 0.00fF
C6434 sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6435 sky130_fd_sc_hd__dfrtn_1_7/a_651_413# VDD 0.00fF
C6436 sky130_fd_sc_hd__dfrtn_1_17/a_193_47# RESET_COUNTERn 0.02fF
C6437 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# DOUT[14] 0.01fF
C6438 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C6439 sky130_fd_sc_hd__dfrtn_1_9/a_543_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C6440 sky130_fd_sc_hd__dfrtn_1_36/a_1270_413# RESET_COUNTERn 0.00fF
C6441 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C6442 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.01fF
C6443 sky130_fd_sc_hd__dfrtp_1_0/a_805_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C6444 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6445 sky130_fd_sc_hd__inv_1_22/A VIN 0.26fF
C6446 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__inv_1_11/Y 0.01fF
C6447 sky130_fd_sc_hd__nor3_2_3/C DOUT[7] 0.13fF
C6448 VDD RESET_COUNTERn 12.19fF
C6449 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C6450 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_761_289# 0.00fF
C6451 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_6/Y 0.02fF
C6452 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_12/A 0.00fF
C6453 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C6454 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C6455 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C6456 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C6457 sky130_fd_sc_hd__or2b_1_0/a_301_297# SEL_CONV_TIME[0] 0.00fF
C6458 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C6459 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C6460 sky130_fd_sc_hd__inv_1_1/Y DOUT[5] 0.00fF
C6461 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6462 sky130_fd_sc_hd__dfrtn_1_27/a_1270_413# DOUT[23] 0.00fF
C6463 sky130_fd_sc_hd__nor3_1_13/a_193_297# sky130_fd_sc_hd__dfrtn_1_10/a_27_47# 0.00fF
C6464 sky130_fd_sc_hd__nor3_1_13/a_109_297# sky130_fd_sc_hd__dfrtn_1_10/a_193_47# 0.00fF
C6465 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# 0.00fF
C6466 CLK_REF sky130_fd_sc_hd__o211a_1_1/a_215_47# 0.00fF
C6467 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C6468 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C6469 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# SEL_CONV_TIME[1] 0.03fF
C6470 sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# 0.00fF
C6471 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_1270_413# 0.00fF
C6472 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_639_47# 0.00fF
C6473 sky130_fd_sc_hd__dfrtn_1_25/a_448_47# sky130_fd_sc_hd__dfrtn_1_27/a_543_47# 0.00fF
C6474 sky130_fd_sc_hd__dfrtn_1_25/a_651_413# sky130_fd_sc_hd__dfrtn_1_27/a_761_289# 0.00fF
C6475 sky130_fd_sc_hd__dfrtn_1_25/a_639_47# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C6476 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_31/a_193_47# 0.00fF
C6477 sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C6478 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C6479 sky130_fd_sc_hd__dfrtn_1_42/a_651_413# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C6480 sky130_fd_sc_hd__nor3_1_4/a_193_297# DOUT[7] 0.00fF
C6481 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__inv_1_33/A 0.02fF
C6482 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_14/a_27_47# 0.01fF
C6483 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C6484 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_12/A 0.03fF
C6485 sky130_fd_sc_hd__dfrtn_1_34/a_805_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C6486 sky130_fd_sc_hd__dfrtn_1_5/a_805_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C6487 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C6488 sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C6489 DOUT[13] sky130_fd_sc_hd__dfrtn_1_34/a_1270_413# 0.00fF
C6490 sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# RESET_COUNTERn 0.02fF
C6491 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# SEL_CONV_TIME[0] 0.03fF
C6492 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__dfrtn_1_33/a_193_47# 0.00fF
C6493 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_33/a_27_47# 0.00fF
C6494 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__dfrtn_1_34/a_651_413# 0.00fF
C6495 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__dfrtn_1_34/a_448_47# 0.00fF
C6496 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__dfrtn_1_14/a_193_47# -0.05fF
C6497 sky130_fd_sc_hd__dfrtn_1_8/a_543_47# sky130_fd_sc_hd__inv_1_9/Y 0.00fF
C6498 sky130_fd_sc_hd__dfrtn_1_28/a_761_289# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C6499 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# CLK_REF 0.00fF
C6500 sky130_fd_sc_hd__dfrtn_1_19/a_651_413# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C6501 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C6502 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__or3b_2_0/a_388_297# 0.00fF
C6503 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__dfrtn_1_22/a_1108_47# -0.00fF
C6504 sky130_fd_sc_hd__dfrtn_1_36/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6505 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C6506 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_23/a_27_47# 0.00fF
C6507 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C6508 sky130_fd_sc_hd__dfrtn_1_27/a_1462_47# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C6509 sky130_fd_sc_hd__a221oi_4_0/a_27_297# SEL_CONV_TIME[3] 0.02fF
C6510 sky130_fd_sc_hd__inv_1_38/Y DOUT[21] 0.25fF
C6511 sky130_fd_sc_hd__or2b_1_0/a_27_53# DOUT[21] 0.00fF
C6512 sky130_fd_sc_hd__dfrtn_1_7/a_639_47# DOUT[14] 0.00fF
C6513 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# VDD 0.05fF
C6514 sky130_fd_sc_hd__dfrtn_1_25/a_1217_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C6515 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# 0.01fF
C6516 sky130_fd_sc_hd__dfrtn_1_39/a_651_413# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C6517 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.03fF
C6518 sky130_fd_sc_hd__dfrtn_1_3/a_761_289# VDD 0.04fF
C6519 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__mux4_2_0/a_1064_47# 0.00fF
C6520 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__inv_1_1/A 0.02fF
C6521 sky130_fd_sc_hd__dfrtn_1_17/a_1462_47# RESET_COUNTERn 0.00fF
C6522 sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C6523 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__o2111a_2_0/a_566_47# -0.00fF
C6524 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# RESET_COUNTERn -0.00fF
C6525 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C6526 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C6527 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C6528 sky130_fd_sc_hd__dfrtn_1_21/a_448_47# sky130_fd_sc_hd__dfrtn_1_19/a_1462_47# 0.00fF
C6529 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_1217_47# 0.00fF
C6530 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C6531 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C6532 DOUT[16] sky130_fd_sc_hd__inv_1_38/A 0.10fF
C6533 sky130_fd_sc_hd__dfrtn_1_36/a_193_47# sky130_fd_sc_hd__inv_1_38/A 0.00fF
C6534 sky130_fd_sc_hd__dfrtn_1_19/a_1283_21# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C6535 sky130_fd_sc_hd__dfrtn_1_0/a_805_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C6536 DOUT[4] sky130_fd_sc_hd__dfrtn_1_35/a_448_47# 0.00fF
C6537 sky130_fd_sc_hd__dfrtn_1_11/a_1217_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C6538 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# 0.00fF
C6539 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_31/a_761_289# 0.00fF
C6540 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C6541 sky130_fd_sc_hd__a221oi_4_0/a_27_297# SEL_CONV_TIME[2] 0.01fF
C6542 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C6543 sky130_fd_sc_hd__dfrtn_1_31/a_805_47# RESET_COUNTERn 0.00fF
C6544 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C6545 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.00fF
C6546 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__dfrtn_1_26/a_761_289# 0.00fF
C6547 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__dfrtn_1_26/a_543_47# 0.00fF
C6548 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C6549 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__dfrtn_1_28/a_27_47# 0.00fF
C6550 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# 0.00fF
C6551 sky130_fd_sc_hd__dfrtn_1_9/a_805_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C6552 sky130_fd_sc_hd__dfrtn_1_32/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6553 sky130_fd_sc_hd__nor3_1_19/Y sky130_fd_sc_hd__nor3_2_3/B 0.23fF
C6554 sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# SEL_CONV_TIME[1] 0.00fF
C6555 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C6556 VDD SEL_CONV_TIME[3] 1.53fF
C6557 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# 0.00fF
C6558 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C6559 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# 0.00fF
C6560 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C6561 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_8/a_1283_21# 0.01fF
C6562 sky130_fd_sc_hd__inv_1_7/Y VDD 0.33fF
C6563 sky130_fd_sc_hd__dfrtn_1_19/a_193_47# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C6564 sky130_fd_sc_hd__dfrtn_1_20/a_639_47# DOUT[2] 0.00fF
C6565 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# sky130_fd_sc_hd__dfrtn_1_16/a_193_47# -0.29fF
C6566 sky130_fd_sc_hd__dfrtn_1_22/a_448_47# sky130_fd_sc_hd__dfrtn_1_23/a_27_47# 0.00fF
C6567 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__dfrtn_1_23/a_448_47# 0.00fF
C6568 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# DOUT[3] 0.00fF
C6569 sky130_fd_sc_hd__dfrtn_1_31/a_1270_413# DONE 0.00fF
C6570 sky130_fd_sc_hd__mux4_2_0/a_1064_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C6571 sky130_fd_sc_hd__o221ai_1_0/a_493_297# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C6572 sky130_fd_sc_hd__dfrtn_1_9/a_651_413# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C6573 sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# sky130_fd_sc_hd__inv_1_27/Y 0.00fF
C6574 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# 0.00fF
C6575 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__dfrtn_1_16/a_27_47# 0.00fF
C6576 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# sky130_fd_sc_hd__inv_1_2/A 0.01fF
C6577 sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# SEL_CONV_TIME[0] 0.00fF
C6578 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_33/a_1217_47# 0.00fF
C6579 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__dfrtn_1_33/a_639_47# 0.00fF
C6580 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__dfrtn_1_33/a_761_289# 0.00fF
C6581 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__dfrtn_1_33/a_651_413# 0.00fF
C6582 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__dfrtn_1_33/a_543_47# 0.00fF
C6583 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__or2_2_0/X 0.01fF
C6584 sky130_fd_sc_hd__dfrtp_1_3/a_1283_21# RESET_COUNTERn 0.03fF
C6585 sky130_fd_sc_hd__o211a_1_0/X RESET_COUNTERn 0.00fF
C6586 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__o211a_1_1/a_215_47# 0.00fF
C6587 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.00fF
C6588 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__o211a_1_1/a_510_47# 0.00fF
C6589 sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C6590 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__nor3_1_19/Y 0.01fF
C6591 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C6592 sky130_fd_sc_hd__dfrtn_1_10/a_639_47# outb 0.00fF
C6593 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C6594 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# DOUT[21] 0.00fF
C6595 sky130_fd_sc_hd__nor3_2_3/B DOUT[14] 2.23fF
C6596 sky130_fd_sc_hd__nor3_1_10/a_193_297# DOUT[14] 0.00fF
C6597 VDD SEL_CONV_TIME[2] 1.82fF
C6598 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_23/a_1217_47# 0.00fF
C6599 sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# VDD 0.09fF
C6600 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6601 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_3/a_761_289# 0.00fF
C6602 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_3/a_27_47# 0.00fF
C6603 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C6604 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__dfrtn_1_3/a_193_47# 0.01fF
C6605 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_543_47# 0.00fF
C6606 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C6607 sky130_fd_sc_hd__dfrtn_1_12/a_805_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C6608 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__inv_1_46/Y 0.00fF
C6609 sky130_fd_sc_hd__dfrtn_1_20/a_543_47# sky130_fd_sc_hd__inv_1_35/Y 0.00fF
C6610 sky130_fd_sc_hd__nor3_1_17/a_193_297# sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# 0.00fF
C6611 sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6612 sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C6613 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__dfrtn_1_38/a_1462_47# 0.00fF
C6614 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# 0.00fF
C6615 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# 0.00fF
C6616 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__dfrtp_1_2/a_761_289# 0.00fF
C6617 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__dfrtp_1_2/a_651_413# 0.00fF
C6618 sky130_fd_sc_hd__dfrtp_1_1/a_448_47# sky130_fd_sc_hd__dfrtp_1_2/a_543_47# 0.00fF
C6619 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# 0.00fF
C6620 sky130_fd_sc_hd__inv_1_10/A RESET_COUNTERn 2.08fF
C6621 sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C6622 sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# RESET_COUNTERn 0.00fF
C6623 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C6624 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# 0.00fF
C6625 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C6626 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C6627 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C6628 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# 0.00fF
C6629 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C6630 sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C6631 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C6632 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# sky130_fd_sc_hd__inv_1_44/Y 0.02fF
C6633 sky130_fd_sc_hd__dfrtn_1_42/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C6634 sky130_fd_sc_hd__dfrtn_1_42/a_1108_47# VDD 0.06fF
C6635 sky130_fd_sc_hd__dfrtn_1_36/a_1462_47# sky130_fd_sc_hd__inv_1_38/A 0.00fF
C6636 sky130_fd_sc_hd__nor3_1_16/a_193_297# VDD 0.00fF
C6637 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# DOUT[14] 0.00fF
C6638 sky130_fd_sc_hd__dfrtn_1_29/a_805_47# DOUT[21] 0.00fF
C6639 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# RESET_COUNTERn 0.02fF
C6640 sky130_fd_sc_hd__or2_2_0/a_121_297# sky130_fd_sc_hd__o211a_1_1/X 0.00fF
C6641 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_25/a_27_47# 0.00fF
C6642 sky130_fd_sc_hd__dfrtn_1_10/a_1283_21# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C6643 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.02fF
C6644 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.02fF
C6645 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# 0.01fF
C6646 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__dfrtn_1_23/a_651_413# -0.00fF
C6647 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# sky130_fd_sc_hd__dfrtn_1_23/a_448_47# -0.00fF
C6648 VDD HEADER_0/a_508_138# 0.05fF
C6649 sky130_fd_sc_hd__inv_1_54/A SEL_CONV_TIME[1] 0.01fF
C6650 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C6651 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# VDD 0.00fF
C6652 SEL_CONV_TIME[1] sky130_fd_sc_hd__inv_1_48/A 0.55fF
C6653 sky130_fd_sc_hd__inv_1_41/Y sky130_fd_sc_hd__inv_1_44/A 0.00fF
C6654 SEL_CONV_TIME[0] sky130_fd_sc_hd__inv_1_48/Y 0.01fF
C6655 sky130_fd_sc_hd__dfrtn_1_9/a_639_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C6656 sky130_fd_sc_hd__dfrtn_1_4/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6657 sky130_fd_sc_hd__dfrtn_1_14/a_651_413# DOUT[11] 0.00fF
C6658 sky130_fd_sc_hd__dfrtn_1_4/a_639_47# VDD 0.00fF
C6659 sky130_fd_sc_hd__dfrtn_1_38/a_651_413# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C6660 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C6661 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# 0.00fF
C6662 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# 0.00fF
C6663 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.02fF
C6664 sky130_fd_sc_hd__dfrtn_1_7/a_651_413# DOUT[3] 0.00fF
C6665 sky130_fd_sc_hd__nor3_1_9/a_193_297# DOUT[14] 0.00fF
C6666 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_29/a_651_413# 0.00fF
C6667 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C6668 sky130_fd_sc_hd__dfrtn_1_19/a_27_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C6669 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.01fF
C6670 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__or2_2_0/a_121_297# 0.00fF
C6671 SLC_0/a_264_22# VDD 0.10fF
C6672 sky130_fd_sc_hd__dfrtp_1_3/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6673 sky130_fd_sc_hd__inv_1_26/A sky130_fd_sc_hd__nor3_2_3/C 0.56fF
C6674 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C6675 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__inv_1_43/A 0.02fF
C6676 sky130_fd_sc_hd__dfrtn_1_16/a_193_47# DOUT[15] 0.01fF
C6677 sky130_fd_sc_hd__dfrtn_1_7/a_651_413# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C6678 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# DOUT[21] 0.00fF
C6679 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__nor3_1_2/a_193_297# 0.00fF
C6680 RESET_COUNTERn DOUT[3] 0.35fF
C6681 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C6682 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.00fF
C6683 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C6684 sky130_fd_sc_hd__nand3b_1_0/a_232_47# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C6685 sky130_fd_sc_hd__dfrtn_1_29/a_805_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C6686 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# sky130_fd_sc_hd__dfrtn_1_7/a_193_47# 0.01fF
C6687 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__dfrtn_1_7/a_27_47# 0.01fF
C6688 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__dfrtn_1_7/a_761_289# 0.01fF
C6689 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# 0.01fF
C6690 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# sky130_fd_sc_hd__dfrtn_1_7/a_543_47# 0.01fF
C6691 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# 0.01fF
C6692 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C6693 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__inv_1_0/Y 0.32fF
C6694 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_0/a_1270_413# 0.00fF
C6695 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_3/a_651_413# 0.00fF
C6696 sky130_fd_sc_hd__nor3_2_2/a_27_297# DOUT[15] 0.02fF
C6697 DOUT[4] sky130_fd_sc_hd__dfrtn_1_12/a_193_47# 0.00fF
C6698 sky130_fd_sc_hd__mux4_2_0/a_1060_369# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C6699 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__dfrtn_1_28/a_639_47# -0.00fF
C6700 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# VDD 0.01fF
C6701 sky130_fd_sc_hd__dfrtp_1_0/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6702 sky130_fd_sc_hd__dfrtn_1_36/a_543_47# sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C6703 sky130_fd_sc_hd__inv_1_2/A RESET_COUNTERn 1.05fF
C6704 VDD DOUT[10] 0.33fF
C6705 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# 0.00fF
C6706 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# 0.00fF
C6707 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__dfrtn_1_6/a_805_47# -0.00fF
C6708 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# -0.00fF
C6709 DOUT[5] RESET_COUNTERn 0.00fF
C6710 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# DOUT[7] 0.01fF
C6711 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# DOUT[6] 0.00fF
C6712 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# DOUT[20] 0.01fF
C6713 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C6714 sky130_fd_sc_hd__dfrtn_1_22/a_448_47# RESET_COUNTERn 0.00fF
C6715 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C6716 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_639_47# 0.00fF
C6717 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C6718 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_805_47# 0.00fF
C6719 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C6720 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C6721 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C6722 sky130_fd_sc_hd__dfrtn_1_39/a_1270_413# VDD 0.00fF
C6723 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__inv_1_50/Y 0.01fF
C6724 CLK_REF sky130_fd_sc_hd__dfrtn_1_20/a_543_47# 0.00fF
C6725 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_32/a_193_47# 0.02fF
C6726 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6727 DOUT[4] sky130_fd_sc_hd__or2b_1_0/X 0.01fF
C6728 sky130_fd_sc_hd__dfrtn_1_30/a_543_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C6729 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_3/a_761_289# 0.00fF
C6730 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_10/a_543_47# -0.00fF
C6731 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# sky130_fd_sc_hd__dfrtn_1_3/a_543_47# 0.00fF
C6732 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__dfrtn_1_3/a_651_413# 0.00fF
C6733 sky130_fd_sc_hd__dfrtn_1_14/a_543_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C6734 sky130_fd_sc_hd__inv_1_14/A sky130_fd_sc_hd__nor3_2_3/C 0.06fF
C6735 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# outb 0.00fF
C6736 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C6737 DOUT[19] sky130_fd_sc_hd__nor3_1_4/A 0.01fF
C6738 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C6739 sky130_fd_sc_hd__dfrtn_1_18/a_1270_413# VDD 0.00fF
C6740 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C6741 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C6742 sky130_fd_sc_hd__dfrtn_1_21/a_448_47# sky130_fd_sc_hd__inv_1_35/Y 0.01fF
C6743 sky130_fd_sc_hd__dfrtn_1_41/a_805_47# DOUT[2] 0.00fF
C6744 sky130_fd_sc_hd__dfrtn_1_21/a_543_47# sky130_fd_sc_hd__inv_1_35/A 0.01fF
C6745 sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.01fF
C6746 sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C6747 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__inv_1_43/A 0.01fF
C6748 sky130_fd_sc_hd__dfrtn_1_16/a_1283_21# RESET_COUNTERn 0.00fF
C6749 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# DOUT[14] 0.00fF
C6750 sky130_fd_sc_hd__dfrtn_1_8/a_1108_47# DOUT[21] 0.00fF
C6751 sky130_fd_sc_hd__dfrtn_1_8/a_27_47# RESET_COUNTERn 0.03fF
C6752 sky130_fd_sc_hd__dfrtn_1_9/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6753 VDD sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.06fF
C6754 sky130_fd_sc_hd__dfrtn_1_20/a_761_289# sky130_fd_sc_hd__dfrtn_1_20/a_543_47# -0.00fF
C6755 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# -0.00fF
C6756 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# -0.00fF
C6757 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_805_47# 0.00fF
C6758 sky130_fd_sc_hd__o211a_1_1/a_297_297# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C6759 sky130_fd_sc_hd__dfrtn_1_41/a_639_47# sky130_fd_sc_hd__dfrtn_1_38/a_543_47# 0.00fF
C6760 sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C6761 sky130_fd_sc_hd__dfrtn_1_41/a_448_47# sky130_fd_sc_hd__dfrtn_1_38/a_448_47# 0.00fF
C6762 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__dfrtn_1_38/a_1270_413# 0.00fF
C6763 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# sky130_fd_sc_hd__dfrtn_1_38/a_805_47# 0.00fF
C6764 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# sky130_fd_sc_hd__dfrtn_1_38/a_639_47# 0.00fF
C6765 sky130_fd_sc_hd__dfrtn_1_19/a_1283_21# VDD 0.09fF
C6766 sky130_fd_sc_hd__dfrtp_1_3/a_651_413# DOUT[23] 0.00fF
C6767 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__conb_1_0/LO 0.00fF
C6768 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__dfrtn_1_1/a_193_47# 0.00fF
C6769 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__dfrtn_1_1/a_27_47# 0.00fF
C6770 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_1/a_543_47# 0.00fF
C6771 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_1/a_805_47# 0.00fF
C6772 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_1/a_651_413# 0.00fF
C6773 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_1/a_639_47# 0.00fF
C6774 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_13/Y 0.07fF
C6775 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_13/A 0.00fF
C6776 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C6777 sky130_fd_sc_hd__o221ai_1_0/a_213_123# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6778 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__mux4_2_0/a_1064_47# 0.00fF
C6779 sky130_fd_sc_hd__nor3_1_17/a_109_297# VDD 0.00fF
C6780 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C6781 sky130_fd_sc_hd__mux4_2_0/a_1279_413# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C6782 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# SEL_CONV_TIME[1] 0.00fF
C6783 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_805_47# -0.00fF
C6784 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C6785 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.06fF
C6786 DONE SEL_CONV_TIME[0] 0.00fF
C6787 sky130_fd_sc_hd__inv_1_35/A sky130_fd_sc_hd__inv_1_35/Y 0.03fF
C6788 sky130_fd_sc_hd__dfrtn_1_33/a_1217_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C6789 sky130_fd_sc_hd__dfrtn_1_16/a_1462_47# DOUT[15] 0.00fF
C6790 DOUT[4] sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C6791 DOUT[4] DOUT[16] 0.02fF
C6792 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C6793 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C6794 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C6795 sky130_fd_sc_hd__dfrtn_1_23/a_1462_47# DOUT[21] 0.00fF
C6796 sky130_fd_sc_hd__dfrtn_1_23/a_651_413# RESET_COUNTERn 0.00fF
C6797 sky130_fd_sc_hd__dfrtn_1_22/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C6798 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__or3b_2_0/a_472_297# 0.00fF
C6799 sky130_fd_sc_hd__nor3_1_1/a_193_297# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C6800 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__dfrtn_1_26/a_639_47# 0.00fF
C6801 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__dfrtn_1_26/a_805_47# 0.00fF
C6802 sky130_fd_sc_hd__dfrtn_1_12/a_1462_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C6803 sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# DOUT[7] 0.00fF
C6804 sky130_fd_sc_hd__dfrtn_1_7/a_543_47# RESET_COUNTERn 0.01fF
C6805 sky130_fd_sc_hd__dfrtn_1_7/a_651_413# DOUT[20] 0.00fF
C6806 sky130_fd_sc_hd__dfrtn_1_7/a_448_47# DOUT[6] 0.00fF
C6807 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_29/a_761_289# 0.00fF
C6808 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C6809 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__mux4_1_0/X 0.01fF
C6810 VDD sky130_fd_sc_hd__or3_1_0/X 0.25fF
C6811 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.00fF
C6812 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__nor3_2_0/A 0.01fF
C6813 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_0/a_448_47# -0.00fF
C6814 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# -0.00fF
C6815 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# RESET_COUNTERn 0.00fF
C6816 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# DOUT[7] 0.00fF
C6817 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# DOUT[6] 0.00fF
C6818 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# CLK_REF 0.02fF
C6819 DOUT[6] DOUT[8] 0.05fF
C6820 DOUT[20] RESET_COUNTERn 1.03fF
C6821 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C6822 sky130_fd_sc_hd__inv_1_7/Y DOUT[3] 0.01fF
C6823 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# DOUT[17] 0.00fF
C6824 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_757_363# -0.00fF
C6825 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__mux4_1_0/a_750_97# -0.00fF
C6826 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_32/a_1462_47# 0.00fF
C6827 sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# sky130_fd_sc_hd__dfrtn_1_27/a_761_289# 0.00fF
C6828 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# sky130_fd_sc_hd__dfrtn_1_27/a_543_47# 0.00fF
C6829 sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C6830 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_448_47# 0.00fF
C6831 sky130_fd_sc_hd__dfrtn_1_26/a_651_413# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C6832 sky130_fd_sc_hd__dfrtn_1_24/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6833 sky130_fd_sc_hd__o2111a_2_0/a_458_47# sky130_fd_sc_hd__o311a_1_0/a_266_47# 0.00fF
C6834 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__inv_1_32/A 0.01fF
C6835 sky130_fd_sc_hd__dfrtn_1_24/a_1270_413# VDD 0.00fF
C6836 sky130_fd_sc_hd__dfrtn_1_16/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6837 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# VDD 0.04fF
C6838 CLK_REF sky130_fd_sc_hd__dfrtn_1_21/a_448_47# 0.00fF
C6839 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6840 sky130_fd_sc_hd__dfrtn_1_11/a_1217_47# outb 0.00fF
C6841 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__inv_1_2/A 0.02fF
C6842 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# SEL_CONV_TIME[0] 0.00fF
C6843 SEL_CONV_TIME[0] sky130_fd_sc_hd__nor3_2_3/B 0.63fF
C6844 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__inv_1_53/A 0.03fF
C6845 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C6846 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_31/a_543_47# 0.00fF
C6847 sky130_fd_sc_hd__nor3_2_2/a_281_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6848 sky130_fd_sc_hd__dfrtn_1_9/a_651_413# DOUT[14] 0.00fF
C6849 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__nor3_1_16/a_193_297# 0.00fF
C6850 sky130_fd_sc_hd__dfrtn_1_33/a_543_47# SEL_CONV_TIME[1] 0.00fF
C6851 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__or2_2_0/A 0.01fF
C6852 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.02fF
C6853 sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C6854 sky130_fd_sc_hd__dfrtn_1_8/a_1217_47# RESET_COUNTERn 0.00fF
C6855 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__or3b_2_0/X 0.01fF
C6856 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_14/a_27_47# 0.00fF
C6857 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# sky130_fd_sc_hd__o211a_1_0/X 0.00fF
C6858 sky130_fd_sc_hd__dfrtn_1_30/a_1270_413# SEL_CONV_TIME[1] 0.00fF
C6859 DOUT[12] VIN 3.26fF
C6860 sky130_fd_sc_hd__dfrtn_1_20/a_639_47# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C6861 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_21/a_27_47# 0.00fF
C6862 sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6863 DOUT[4] sky130_fd_sc_hd__or3b_2_0/a_472_297# 0.00fF
C6864 sky130_fd_sc_hd__nand3b_1_1/Y sky130_fd_sc_hd__inv_1_42/A 0.00fF
C6865 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# 0.00fF
C6866 sky130_fd_sc_hd__or3b_2_0/a_388_297# sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# 0.00fF
C6867 VDD sky130_fd_sc_hd__nor3_2_2/A 0.55fF
C6868 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C6869 sky130_fd_sc_hd__dfrtn_1_24/a_805_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C6870 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.00fF
C6871 CLK_REF sky130_fd_sc_hd__inv_1_35/A 0.01fF
C6872 sky130_fd_sc_hd__or3_1_0/a_183_297# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C6873 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6874 sky130_fd_sc_hd__nand3b_1_1/a_53_93# SEL_CONV_TIME[0] 0.02fF
C6875 sky130_fd_sc_hd__or3_1_0/a_29_53# SEL_CONV_TIME[0] 0.01fF
C6876 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C6877 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__nor3_1_3/a_193_297# 0.00fF
C6878 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C6879 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# VDD 0.05fF
C6880 sky130_fd_sc_hd__dfrtn_1_42/a_193_47# sky130_fd_sc_hd__dfrtn_1_23/a_27_47# 0.00fF
C6881 sky130_fd_sc_hd__dfrtn_1_38/a_193_47# SEL_CONV_TIME[1] 0.00fF
C6882 DOUT[4] sky130_fd_sc_hd__dfrtn_1_36/a_1462_47# 0.00fF
C6883 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C6884 sky130_fd_sc_hd__dfrtn_1_34/a_805_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C6885 sky130_fd_sc_hd__or3b_2_0/X sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C6886 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__dfrtn_1_30/a_27_47# 0.00fF
C6887 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__inv_1_36/Y 0.02fF
C6888 sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C6889 VDD sky130_fd_sc_hd__inv_1_53/A 1.03fF
C6890 sky130_fd_sc_hd__dfrtn_1_33/a_761_289# VDD 0.04fF
C6891 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.03fF
C6892 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__o2111a_2_0/X 0.01fF
C6893 sky130_fd_sc_hd__o311a_1_0/a_266_47# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C6894 HEADER_0/a_508_138# DOUT[3] 0.01fF
C6895 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# sky130_fd_sc_hd__inv_1_40/Y 0.00fF
C6896 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__inv_1_27/Y 0.02fF
C6897 sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6898 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C6899 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# DOUT[3] 0.00fF
C6900 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__nand2_1_1/a_113_47# 0.00fF
C6901 sky130_fd_sc_hd__dfrtn_1_30/a_651_413# VDD 0.01fF
C6902 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C6903 sky130_fd_sc_hd__dfrtn_1_4/a_639_47# DOUT[3] 0.00fF
C6904 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__a221oi_4_0/a_1241_47# 0.00fF
C6905 sky130_fd_sc_hd__dfrtn_1_20/a_761_289# sky130_fd_sc_hd__inv_1_35/A 0.02fF
C6906 sky130_fd_sc_hd__dfrtn_1_16/a_651_413# DOUT[23] 0.00fF
C6907 DOUT[4] sky130_fd_sc_hd__dfrtn_1_31/a_543_47# 0.00fF
C6908 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__inv_1_41/Y 0.01fF
C6909 sky130_fd_sc_hd__dfrtn_1_30/a_448_47# sky130_fd_sc_hd__dfrtn_1_31/a_27_47# 0.00fF
C6910 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_448_47# 0.00fF
C6911 sky130_fd_sc_hd__inv_1_2/A HEADER_0/a_508_138# 0.00fF
C6912 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C6913 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# DOUT[14] 0.00fF
C6914 sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C6915 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C6916 sky130_fd_sc_hd__dfrtn_1_4/a_639_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C6917 sky130_fd_sc_hd__dfrtn_1_20/a_1462_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C6918 sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# DOUT[17] 0.00fF
C6919 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_834_97# -0.00fF
C6920 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C6921 sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# sky130_fd_sc_hd__dfrtn_1_27/a_448_47# 0.00fF
C6922 sky130_fd_sc_hd__inv_1_3/A VIN 0.11fF
C6923 sky130_fd_sc_hd__o211a_1_1/a_510_47# sky130_fd_sc_hd__dfrtn_1_17/a_761_289# 0.00fF
C6924 sky130_fd_sc_hd__o211a_1_1/a_215_47# sky130_fd_sc_hd__dfrtn_1_17/a_543_47# 0.00fF
C6925 sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# SEL_CONV_TIME[1] 0.01fF
C6926 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C6927 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_761_289# 0.00fF
C6928 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C6929 sky130_fd_sc_hd__dfrtn_1_25/a_448_47# SEL_CONV_TIME[0] 0.00fF
C6930 sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__o211a_1_0/a_215_47# 0.01fF
C6931 sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6932 sky130_fd_sc_hd__nor3_1_7/a_109_297# DOUT[19] 0.00fF
C6933 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# VDD 0.26fF
C6934 sky130_fd_sc_hd__dfrtn_1_36/a_639_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C6935 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C6936 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# 0.00fF
C6937 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__dfrtn_1_11/a_543_47# 0.00fF
C6938 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_448_47# 0.00fF
C6939 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__dfrtn_1_11/a_27_47# 0.00fF
C6940 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# 0.00fF
C6941 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C6942 sky130_fd_sc_hd__o211a_1_1/a_215_47# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C6943 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__inv_1_22/Y 0.04fF
C6944 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C6945 sky130_fd_sc_hd__inv_1_7/Y DOUT[20] 0.14fF
C6946 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_12/a_805_47# 0.00fF
C6947 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# 0.00fF
C6948 DOUT[4] sky130_fd_sc_hd__dfrtn_1_32/a_1270_413# 0.00fF
C6949 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C6950 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/a_761_289# -0.00fF
C6951 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_1/a_543_47# -0.00fF
C6952 sky130_fd_sc_hd__dfrtn_1_12/a_651_413# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C6953 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# sky130_fd_sc_hd__inv_1_6/A 0.02fF
C6954 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# 0.00fF
C6955 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# 0.00fF
C6956 sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C6957 sky130_fd_sc_hd__dfrtp_1_2/a_805_47# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C6958 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_17/a_639_47# 0.00fF
C6959 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_805_47# 0.00fF
C6960 sky130_fd_sc_hd__nand2_1_1/Y SEL_CONV_TIME[0] 0.00fF
C6961 sky130_fd_sc_hd__inv_1_28/A sky130_fd_sc_hd__or2_2_0/A 0.00fF
C6962 sky130_fd_sc_hd__inv_1_2/A DOUT[10] 0.01fF
C6963 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# 0.00fF
C6964 sky130_fd_sc_hd__dfrtn_1_12/a_651_413# sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# 0.00fF
C6965 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_14/a_805_47# 0.00fF
C6966 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# 0.00fF
C6967 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# 0.00fF
C6968 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_37/a_761_289# -0.00fF
C6969 VDD sky130_fd_sc_hd__inv_1_4/Y 0.24fF
C6970 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C6971 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# 0.00fF
C6972 sky130_fd_sc_hd__dfrtn_1_28/a_543_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C6973 sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__or2_2_0/B 0.44fF
C6974 sky130_fd_sc_hd__inv_1_42/Y VDD 0.42fF
C6975 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6976 sky130_fd_sc_hd__dfrtn_1_26/a_761_289# VDD 0.05fF
C6977 sky130_fd_sc_hd__o211a_1_0/a_215_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C6978 sky130_fd_sc_hd__nor3_2_3/C VIN 0.08fF
C6979 CLK_REF sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C6980 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C6981 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# DOUT[14] 0.02fF
C6982 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6983 sky130_fd_sc_hd__nor3_2_0/a_27_297# sky130_fd_sc_hd__nor3_2_3/B 0.03fF
C6984 DOUT[4] sky130_fd_sc_hd__or2b_1_0/a_219_297# 0.00fF
C6985 sky130_fd_sc_hd__dfrtn_1_34/a_543_47# VDD 0.06fF
C6986 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_7/a_27_47# 0.00fF
C6987 sky130_fd_sc_hd__dfrtp_1_2/a_805_47# VDD 0.00fF
C6988 DOUT[9] DOUT[18] 0.02fF
C6989 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__dfrtn_1_30/a_543_47# 0.00fF
C6990 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__dfrtn_1_30/a_761_289# 0.00fF
C6991 sky130_fd_sc_hd__dfrtn_1_23/a_761_289# sky130_fd_sc_hd__inv_1_40/Y 0.02fF
C6992 sky130_fd_sc_hd__dfrtn_1_28/a_543_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C6993 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C6994 sky130_fd_sc_hd__dfrtn_1_16/a_448_47# sky130_fd_sc_hd__inv_1_26/A 0.00fF
C6995 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C6996 sky130_fd_sc_hd__o2111a_2_0/a_80_21# SEL_CONV_TIME[1] 0.02fF
C6997 sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# DOUT[21] 0.01fF
C6998 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# RESET_COUNTERn 0.01fF
C6999 sky130_fd_sc_hd__dfrtn_1_12/a_805_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C7000 sky130_fd_sc_hd__dfrtn_1_42/a_1462_47# sky130_fd_sc_hd__dfrtn_1_23/a_27_47# 0.00fF
C7001 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_6/a_448_47# 0.00fF
C7002 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C7003 sky130_fd_sc_hd__dfrtn_1_37/a_805_47# RESET_COUNTERn 0.00fF
C7004 sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# sky130_fd_sc_hd__inv_1_36/A 0.01fF
C7005 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_13/Y 0.02fF
C7006 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C7007 DOUT[9] sky130_fd_sc_hd__dfrtn_1_6/a_543_47# 0.00fF
C7008 sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# DOUT[3] 0.00fF
C7009 DOUT[13] SEL_CONV_TIME[1] 0.24fF
C7010 sky130_fd_sc_hd__nor3_1_4/a_193_297# VIN 0.00fF
C7011 sky130_fd_sc_hd__dfrtn_1_33/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7012 sky130_fd_sc_hd__dfrtn_1_3/a_639_47# RESET_COUNTERn 0.00fF
C7013 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# DOUT[15] 0.00fF
C7014 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__inv_1_49/A 0.01fF
C7015 sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C7016 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C7017 sky130_fd_sc_hd__dfrtn_1_7/a_543_47# HEADER_0/a_508_138# 0.00fF
C7018 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C7019 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# VDD 0.01fF
C7020 sky130_fd_sc_hd__dfrtn_1_42/a_193_47# RESET_COUNTERn 0.01fF
C7021 sky130_fd_sc_hd__dfrtn_1_21/a_639_47# sky130_fd_sc_hd__inv_1_35/A 0.00fF
C7022 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_10/a_193_47# 0.10fF
C7023 sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# sky130_fd_sc_hd__inv_1_15/A 0.02fF
C7024 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C7025 sky130_fd_sc_hd__nor3_1_5/A DOUT[11] 0.05fF
C7026 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtp_1_3/a_543_47# 0.00fF
C7027 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C7028 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C7029 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C7030 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C7031 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# HEADER_0/a_508_138# 0.00fF
C7032 sky130_fd_sc_hd__dfrtn_1_0/a_1270_413# DOUT[17] 0.00fF
C7033 HEADER_0/a_508_138# DOUT[20] 0.01fF
C7034 sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C7035 sky130_fd_sc_hd__inv_1_38/A RESET_COUNTERn 0.05fF
C7036 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# DOUT[20] 0.00fF
C7037 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# RESET_COUNTERn 0.02fF
C7038 sky130_fd_sc_hd__dfrtn_1_24/a_805_47# sky130_fd_sc_hd__dfrtn_1_29/a_543_47# 0.00fF
C7039 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# sky130_fd_sc_hd__dfrtn_1_29/a_805_47# 0.00fF
C7040 sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# RESET_COUNTERn 0.01fF
C7041 sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# VDD 0.00fF
C7042 sky130_fd_sc_hd__dfrtn_1_33/a_639_47# sky130_fd_sc_hd__inv_1_45/A 0.00fF
C7043 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_34/a_1462_47# 0.00fF
C7044 sky130_fd_sc_hd__dfrtn_1_21/a_193_47# RESET_COUNTERn 0.06fF
C7045 sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# sky130_fd_sc_hd__dfrtn_1_11/a_1462_47# 0.00fF
C7046 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__dfrtn_1_11/a_1217_47# 0.00fF
C7047 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__inv_1_49/A 0.26fF
C7048 sky130_fd_sc_hd__dfrtn_1_42/a_639_47# DOUT[15] 0.00fF
C7049 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7050 sky130_fd_sc_hd__nor3_2_0/A sky130_fd_sc_hd__inv_1_13/A 0.01fF
C7051 DOUT[23] sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C7052 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C7053 sky130_fd_sc_hd__dfrtn_1_14/a_543_47# VDD 0.06fF
C7054 sky130_fd_sc_hd__dfrtn_1_12/a_1270_413# sky130_fd_sc_hd__dfrtn_1_0/a_27_47# 0.00fF
C7055 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__dfrtn_1_34/a_651_413# 0.00fF
C7056 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_0/a_1270_413# 0.00fF
C7057 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# 0.00fF
C7058 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# sky130_fd_sc_hd__dfrtn_1_0/a_543_47# 0.00fF
C7059 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# 0.00fF
C7060 sky130_fd_sc_hd__inv_1_32/A sky130_fd_sc_hd__inv_1_53/Y 0.01fF
C7061 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_0/a_761_289# 0.00fF
C7062 sky130_fd_sc_hd__dfrtn_1_37/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7063 sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7064 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# DOUT[3] 0.00fF
C7065 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# RESET_COUNTERn 0.01fF
C7066 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C7067 sky130_fd_sc_hd__dfrtn_1_34/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7068 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_41/a_651_413# -0.00fF
C7069 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__dfrtn_1_41/a_448_47# -0.00fF
C7070 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C7071 sky130_fd_sc_hd__dfrtn_1_3/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7072 sky130_fd_sc_hd__inv_1_48/A DOUT[21] 0.13fF
C7073 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_8/a_1270_413# 0.00fF
C7074 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# lc_out 0.01fF
C7075 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C7076 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# -0.00fF
C7077 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__inv_1_2/A 0.01fF
C7078 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__nor3_1_5/a_109_297# 0.00fF
C7079 sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# RESET_COUNTERn 0.03fF
C7080 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__inv_1_51/Y 0.01fF
C7081 sky130_fd_sc_hd__dfrtn_1_22/a_761_289# sky130_fd_sc_hd__inv_1_39/Y 0.02fF
C7082 sky130_fd_sc_hd__dfrtn_1_25/a_1217_47# RESET_COUNTERn 0.00fF
C7083 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__nor3_2_3/C 1.31fF
C7084 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C7085 sky130_fd_sc_hd__dfrtp_1_3/a_651_413# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C7086 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# sky130_fd_sc_hd__inv_1_32/Y 0.00fF
C7087 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C7088 sky130_fd_sc_hd__inv_1_11/Y RESET_COUNTERn 0.68fF
C7089 sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# RESET_COUNTERn 0.02fF
C7090 sky130_fd_sc_hd__dfrtp_1_0/a_1217_47# DOUT[15] 0.00fF
C7091 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_26/a_639_47# 0.00fF
C7092 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.05fF
C7093 sky130_fd_sc_hd__nor3_1_10/a_193_297# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C7094 sky130_fd_sc_hd__or2_2_0/a_39_297# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C7095 sky130_fd_sc_hd__dfrtn_1_4/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7096 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# SEL_CONV_TIME[3] 0.00fF
C7097 en DOUT[7] 0.03fF
C7098 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_651_413# 0.00fF
C7099 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C7100 sky130_fd_sc_hd__dfrtn_1_28/a_1270_413# SEL_CONV_TIME[1] 0.00fF
C7101 sky130_fd_sc_hd__inv_1_44/A sky130_fd_sc_hd__or3_1_0/C 0.00fF
C7102 sky130_fd_sc_hd__o311a_1_0/A3 sky130_fd_sc_hd__inv_1_48/A 0.01fF
C7103 sky130_fd_sc_hd__mux4_2_0/a_1281_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C7104 sky130_fd_sc_hd__dfrtn_1_42/a_1462_47# RESET_COUNTERn 0.00fF
C7105 sky130_fd_sc_hd__dfrtn_1_37/a_805_47# SEL_CONV_TIME[3] 0.00fF
C7106 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# DOUT[3] 0.00fF
C7107 DOUT[9] DOUT[22] 0.30fF
C7108 sky130_fd_sc_hd__mux4_2_0/a_1279_413# sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.00fF
C7109 sky130_fd_sc_hd__inv_1_3/Y RESET_COUNTERn 0.47fF
C7110 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# RESET_COUNTERn 0.02fF
C7111 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_10/a_1462_47# 0.00fF
C7112 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtp_1_3/a_805_47# 0.00fF
C7113 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtp_1_3/a_639_47# 0.00fF
C7114 sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# sky130_fd_sc_hd__dfrtp_1_3/a_761_289# 0.00fF
C7115 sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# sky130_fd_sc_hd__dfrtp_1_3/a_543_47# 0.00fF
C7116 sky130_fd_sc_hd__or2b_1_0/X sky130_fd_sc_hd__inv_1_44/A 0.01fF
C7117 sky130_fd_sc_hd__dfrtn_1_19/a_27_47# RESET_COUNTERn 0.04fF
C7118 CLK_REF sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# 0.01fF
C7119 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__inv_1_2/A 0.01fF
C7120 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__inv_1_43/A 0.01fF
C7121 sky130_fd_sc_hd__dfrtn_1_24/a_1462_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C7122 sky130_fd_sc_hd__mux4_2_0/a_193_369# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C7123 sky130_fd_sc_hd__dfrtn_1_24/a_805_47# SEL_CONV_TIME[0] 0.00fF
C7124 sky130_fd_sc_hd__inv_1_29/Y RESET_COUNTERn 0.00fF
C7125 sky130_fd_sc_hd__o221ai_1_0/a_493_297# RESET_COUNTERn 0.00fF
C7126 sky130_fd_sc_hd__nor3_1_17/a_193_297# DOUT[21] 0.00fF
C7127 sky130_fd_sc_hd__or3_1_0/a_111_297# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C7128 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__o2111a_2_0/a_386_47# 0.00fF
C7129 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C7130 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C7131 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__inv_1_8/A 0.34fF
C7132 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_543_47# -0.00fF
C7133 sky130_fd_sc_hd__nor3_2_1/a_27_297# sky130_fd_sc_hd__conb_1_0/LO 0.00fF
C7134 sky130_fd_sc_hd__dfrtn_1_31/a_1217_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C7135 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.00fF
C7136 sky130_fd_sc_hd__dfrtn_1_35/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_543_47# 0.00fF
C7137 sky130_fd_sc_hd__dfrtn_1_35/a_543_47# sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C7138 DOUT[13] sky130_fd_sc_hd__dfrtn_1_31/a_639_47# 0.00fF
C7139 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.01fF
C7140 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# 0.00fF
C7141 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# sky130_fd_sc_hd__dfrtn_1_39/a_193_47# 0.00fF
C7142 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_651_413# 0.00fF
C7143 sky130_fd_sc_hd__dfrtn_1_37/a_805_47# SEL_CONV_TIME[2] 0.00fF
C7144 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_29/a_639_47# 0.00fF
C7145 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C7146 sky130_fd_sc_hd__dfrtn_1_28/a_651_413# VDD 0.01fF
C7147 sky130_fd_sc_hd__dfrtn_1_23/a_543_47# sky130_fd_sc_hd__inv_1_39/Y 0.00fF
C7148 sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# sky130_fd_sc_hd__inv_1_7/Y 0.01fF
C7149 sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7150 sky130_fd_sc_hd__dfrtn_1_25/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7151 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_37/a_761_289# 0.01fF
C7152 sky130_fd_sc_hd__dfrtn_1_9/a_543_47# sky130_fd_sc_hd__inv_1_12/A 0.02fF
C7153 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# VDD 0.18fF
C7154 sky130_fd_sc_hd__dfrtn_1_16/a_1283_21# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C7155 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__inv_1_50/Y 0.01fF
C7156 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__inv_1_46/Y 0.00fF
C7157 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C7158 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C7159 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__inv_1_14/A 0.02fF
C7160 sky130_fd_sc_hd__mux4_1_0/a_1290_413# SEL_CONV_TIME[1] 0.03fF
C7161 sky130_fd_sc_hd__nor3_1_10/a_109_297# DOUT[9] 0.00fF
C7162 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C7163 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.01fF
C7164 sky130_fd_sc_hd__nor3_1_20/a_193_297# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C7165 DOUT[9] sky130_fd_sc_hd__dfrtn_1_3/a_543_47# 0.00fF
C7166 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__inv_1_40/Y 0.21fF
C7167 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C7168 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_6/A 0.39fF
C7169 VDD sky130_fd_sc_hd__inv_1_47/A 0.32fF
C7170 sky130_fd_sc_hd__dfrtn_1_39/a_193_47# sky130_fd_sc_hd__inv_1_32/Y 0.06fF
C7171 sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# VDD 0.08fF
C7172 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C7173 sky130_fd_sc_hd__dfrtn_1_42/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7174 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# DOUT[21] 0.00fF
C7175 sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# RESET_COUNTERn -0.00fF
C7176 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# DOUT[20] 0.00fF
C7177 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C7178 sky130_fd_sc_hd__inv_1_49/Y RESET_COUNTERn 0.02fF
C7179 sky130_fd_sc_hd__inv_1_11/A sky130_fd_sc_hd__nor3_2_3/C 0.07fF
C7180 sky130_fd_sc_hd__mux4_2_0/a_872_316# sky130_fd_sc_hd__nand2_1_1/a_113_47# 0.00fF
C7181 sky130_fd_sc_hd__inv_1_4/Y DOUT[3] 0.00fF
C7182 sky130_fd_sc_hd__dfrtp_1_3/a_1270_413# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C7183 DOUT[1] sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# 0.00fF
C7184 DOUT[4] sky130_fd_sc_hd__dfrtn_1_8/a_1283_21# 0.00fF
C7185 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_4/a_761_289# 0.00fF
C7186 sky130_fd_sc_hd__dfrtn_1_23/a_651_413# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C7187 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_26/a_448_47# 0.00fF
C7188 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7189 sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# SEL_CONV_TIME[3] 0.00fF
C7190 sky130_fd_sc_hd__dfrtn_1_16/a_761_289# DOUT[2] 0.01fF
C7191 sky130_fd_sc_hd__dfrtn_1_42/a_193_47# sky130_fd_sc_hd__dfrtn_1_42/a_1108_47# -0.00fF
C7192 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# sky130_fd_sc_hd__dfrtn_1_42/a_448_47# -0.00fF
C7193 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_27_47# 0.00fF
C7194 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_4/Y 0.01fF
C7195 sky130_fd_sc_hd__dfrtn_1_30/a_639_47# SEL_CONV_TIME[0] 0.00fF
C7196 sky130_fd_sc_hd__nor3_1_4/a_109_297# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C7197 sky130_fd_sc_hd__mux4_1_0/a_750_97# VDD 0.03fF
C7198 sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7199 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C7200 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C7201 DOUT[15] sky130_fd_sc_hd__inv_1_39/Y 0.00fF
C7202 sky130_fd_sc_hd__dfrtn_1_10/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7203 sky130_fd_sc_hd__dfrtn_1_10/a_805_47# VDD 0.00fF
C7204 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_19/a_543_47# 0.00fF
C7205 sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# RESET_COUNTERn 0.00fF
C7206 sky130_fd_sc_hd__nor3_2_2/a_281_297# DOUT[2] 0.01fF
C7207 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# VIN 0.13fF
C7208 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# sky130_fd_sc_hd__dfrtn_1_15/a_193_47# 0.00fF
C7209 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# 0.00fF
C7210 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# 0.00fF
C7211 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# sky130_fd_sc_hd__dfrtn_1_15/a_761_289# 0.00fF
C7212 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_651_413# 0.00fF
C7213 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# DOUT[23] 0.00fF
C7214 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C7215 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_20/a_193_47# 0.01fF
C7216 sky130_fd_sc_hd__nor3_1_3/a_193_297# DOUT[19] 0.00fF
C7217 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C7218 sky130_fd_sc_hd__nor3_1_16/a_193_297# sky130_fd_sc_hd__inv_1_38/A 0.00fF
C7219 sky130_fd_sc_hd__dfrtn_1_27/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_543_47# -0.00fF
C7220 sky130_fd_sc_hd__nor3_1_9/a_109_297# DOUT[9] 0.00fF
C7221 sky130_fd_sc_hd__dfrtn_1_19/a_1217_47# RESET_COUNTERn 0.00fF
C7222 sky130_fd_sc_hd__nor3_1_8/a_193_297# RESET_COUNTERn 0.00fF
C7223 sky130_fd_sc_hd__inv_1_17/A sky130_fd_sc_hd__inv_1_24/A 0.01fF
C7224 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C7225 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_11/a_543_47# 0.00fF
C7226 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C7227 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C7228 sky130_fd_sc_hd__dfrtn_1_38/a_761_289# SEL_CONV_TIME[0] 0.00fF
C7229 sky130_fd_sc_hd__mux4_2_0/a_872_316# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C7230 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_651_413# -0.00fF
C7231 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# DOUT[20] 0.00fF
C7232 sky130_fd_sc_hd__dfrtp_1_0/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7233 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_4/a_639_47# 0.00fF
C7234 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_4/a_651_413# 0.00fF
C7235 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C7236 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_4/a_448_47# 0.00fF
C7237 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C7238 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__dfrtn_1_4/a_543_47# 0.00fF
C7239 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C7240 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_193_47# -0.00fF
C7241 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__dfrtn_1_29/a_543_47# 0.00fF
C7242 sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# SEL_CONV_TIME[2] 0.01fF
C7243 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C7244 DOUT[9] sky130_fd_sc_hd__inv_1_6/A 0.00fF
C7245 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.00fF
C7246 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__inv_1_45/A 0.27fF
C7247 sky130_fd_sc_hd__inv_1_37/A sky130_fd_sc_hd__inv_1_5/Y 0.01fF
C7248 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.00fF
C7249 sky130_fd_sc_hd__inv_1_36/Y sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C7250 sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# SEL_CONV_TIME[2] 0.00fF
C7251 DOUT[1] sky130_fd_sc_hd__dfrtn_1_32/a_193_47# 0.01fF
C7252 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C7253 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C7254 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.00fF
C7255 sky130_fd_sc_hd__dfrtn_1_12/a_805_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C7256 sky130_fd_sc_hd__dfrtn_1_35/a_651_413# VDD 0.01fF
C7257 sky130_fd_sc_hd__dfrtn_1_0/a_1217_47# VDD 0.00fF
C7258 DOUT[4] RESET_COUNTERn 0.13fF
C7259 sky130_fd_sc_hd__inv_1_0/Y RESET_COUNTERn 0.34fF
C7260 sky130_fd_sc_hd__dfrtn_1_12/a_651_413# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C7261 sky130_fd_sc_hd__o311a_1_0/a_368_297# SEL_CONV_TIME[1] 0.00fF
C7262 sky130_fd_sc_hd__dfrtn_1_30/a_543_47# RESET_COUNTERn 0.01fF
C7263 sky130_fd_sc_hd__nor3_1_13/a_193_297# sky130_fd_sc_hd__dfrtn_1_8/a_448_47# 0.00fF
C7264 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C7265 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C7266 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# SEL_CONV_TIME[0] 0.01fF
C7267 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C7268 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__or3b_2_0/X 0.01fF
C7269 sky130_fd_sc_hd__dfrtn_1_18/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_193_47# -0.03fF
C7270 sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C7271 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# DOUT[19] 0.01fF
C7272 sky130_fd_sc_hd__dfrtn_1_27/a_448_47# sky130_fd_sc_hd__or3_1_0/C 0.02fF
C7273 sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# SEL_CONV_TIME[0] 0.00fF
C7274 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_1_22/A 0.01fF
C7275 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# VDD 0.10fF
C7276 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C7277 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_14/a_805_47# 0.00fF
C7278 sky130_fd_sc_hd__dfrtn_1_23/a_1270_413# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C7279 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C7280 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# 0.01fF
C7281 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_24/a_651_413# 0.00fF
C7282 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C7283 sky130_fd_sc_hd__dfrtn_1_39/a_1462_47# sky130_fd_sc_hd__inv_1_32/Y 0.00fF
C7284 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# DONE 0.00fF
C7285 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_651_413# -0.00fF
C7286 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# SLC_0/a_264_22# 0.00fF
C7287 sky130_fd_sc_hd__dfrtp_1_0/a_761_289# SLC_0/a_919_243# 0.00fF
C7288 sky130_fd_sc_hd__dfrtn_1_5/a_805_47# RESET_COUNTERn 0.00fF
C7289 sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C7290 sky130_fd_sc_hd__dfrtp_1_0/a_1108_47# sky130_fd_sc_hd__inv_1_26/A 0.01fF
C7291 sky130_fd_sc_hd__dfrtn_1_9/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7292 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__nand3b_1_0/a_316_47# 0.00fF
C7293 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__nand3b_1_0/a_53_93# 0.00fF
C7294 sky130_fd_sc_hd__inv_1_39/A sky130_fd_sc_hd__nor3_2_3/C 0.29fF
C7295 sky130_fd_sc_hd__dfrtn_1_18/a_1462_47# sky130_fd_sc_hd__inv_1_32/Y 0.00fF
C7296 CLK_REF sky130_fd_sc_hd__dfrtp_1_3/a_651_413# 0.00fF
C7297 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__dfrtn_1_24/a_761_289# 0.00fF
C7298 sky130_fd_sc_hd__dfrtn_1_17/a_193_47# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C7299 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_2/a_805_47# 0.00fF
C7300 sky130_fd_sc_hd__dfrtn_1_7/a_543_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C7301 sky130_fd_sc_hd__o211a_1_1/a_79_21# RESET_COUNTERn 0.01fF
C7302 sky130_fd_sc_hd__dfrtn_1_8/a_1283_21# outb 0.00fF
C7303 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_12/a_805_47# -0.00fF
C7304 sky130_fd_sc_hd__dfrtn_1_10/a_639_47# sky130_fd_sc_hd__dfrtn_1_13/a_761_289# 0.00fF
C7305 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# 0.00fF
C7306 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# 0.00fF
C7307 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# 0.00fF
C7308 sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# VIN 0.05fF
C7309 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# DOUT[11] 0.00fF
C7310 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__inv_1_5/Y 0.02fF
C7311 sky130_fd_sc_hd__o311a_1_0/a_266_297# VDD 0.00fF
C7312 DOUT[9] sky130_fd_sc_hd__dfrtn_1_4/a_805_47# 0.00fF
C7313 sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# SEL_CONV_TIME[3] 0.00fF
C7314 sky130_fd_sc_hd__inv_1_47/Y RESET_COUNTERn 0.24fF
C7315 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C7316 sky130_fd_sc_hd__mux4_2_0/a_288_47# VDD 0.03fF
C7317 sky130_fd_sc_hd__dfrtp_1_0/a_761_289# out 0.01fF
C7318 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# DOUT[0] 0.00fF
C7319 sky130_fd_sc_hd__or2_2_0/a_39_297# VDD 0.10fF
C7320 sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.00fF
C7321 sky130_fd_sc_hd__inv_1_4/Y DOUT[20] 0.02fF
C7322 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# SEL_CONV_TIME[1] 0.00fF
C7323 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# VIN 0.00fF
C7324 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# 0.00fF
C7325 sky130_fd_sc_hd__dfrtn_1_34/a_651_413# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C7326 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__nor3_2_1/a_27_297# 0.00fF
C7327 VIN DOUT[7] 0.09fF
C7328 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_20/a_1462_47# 0.00fF
C7329 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C7330 sky130_fd_sc_hd__o2111a_2_0/a_458_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C7331 sky130_fd_sc_hd__o2111a_2_0/a_674_297# SEL_CONV_TIME[0] 0.00fF
C7332 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C7333 sky130_fd_sc_hd__dfrtn_1_35/a_761_289# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C7334 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# VDD 0.09fF
C7335 sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C7336 sky130_fd_sc_hd__dfrtp_1_2/a_448_47# RESET_COUNTERn 0.00fF
C7337 sky130_fd_sc_hd__dfrtn_1_35/a_193_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C7338 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C7339 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7340 sky130_fd_sc_hd__dfrtn_1_41/a_448_47# VDD 0.03fF
C7341 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7342 sky130_fd_sc_hd__nor3_1_4/a_109_297# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C7343 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# DOUT[7] 0.00fF
C7344 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# RESET_COUNTERn 0.00fF
C7345 sky130_fd_sc_hd__nand2_1_1/a_113_47# SEL_CONV_TIME[1] 0.00fF
C7346 sky130_fd_sc_hd__dfrtn_1_3/a_761_289# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C7347 sky130_fd_sc_hd__nor3_1_19/a_109_297# SEL_CONV_TIME[0] 0.00fF
C7348 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_34/a_193_47# 0.00fF
C7349 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_2/Y 0.26fF
C7350 sky130_fd_sc_hd__nand3b_1_0/a_232_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7351 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_39/a_651_413# 0.00fF
C7352 sky130_fd_sc_hd__dfrtn_1_21/a_193_47# sky130_fd_sc_hd__dfrtn_1_19/a_1283_21# 0.01fF
C7353 sky130_fd_sc_hd__o311a_1_0/a_266_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C7354 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_1462_47# 0.00fF
C7355 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C7356 sky130_fd_sc_hd__dfrtn_1_33/a_639_47# RESET_COUNTERn 0.00fF
C7357 DOUT[1] sky130_fd_sc_hd__dfrtn_1_32/a_1462_47# 0.00fF
C7358 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__dfrtn_1_14/a_651_413# 0.00fF
C7359 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__dfrtn_1_14/a_448_47# 0.00fF
C7360 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C7361 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__mux4_2_0/a_1281_47# 0.00fF
C7362 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__mux4_2_0/a_1064_47# 0.00fF
C7363 sky130_fd_sc_hd__nor3_2_0/A sky130_fd_sc_hd__nor3_2_3/C 0.08fF
C7364 outb sky130_fd_sc_hd__inv_1_23/A 0.03fF
C7365 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__nor3_1_19/Y 0.01fF
C7366 sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7367 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_18/a_651_413# 0.00fF
C7368 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__inv_1_8/Y -0.02fF
C7369 outb RESET_COUNTERn 0.17fF
C7370 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C7371 sky130_fd_sc_hd__dfrtn_1_3/a_651_413# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C7372 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# 0.00fF
C7373 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# 0.00fF
C7374 sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C7375 sky130_fd_sc_hd__nor3_2_3/C DOUT[17] 0.08fF
C7376 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# RESET_COUNTERn 0.02fF
C7377 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtp_1_1/D 0.00fF
C7378 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C7379 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C7380 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C7381 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# sky130_fd_sc_hd__inv_1_47/A 0.01fF
C7382 sky130_fd_sc_hd__o2111a_2_0/a_80_21# DOUT[21] 0.00fF
C7383 SEL_CONV_TIME[1] sky130_fd_sc_hd__inv_1_44/Y 0.14fF
C7384 sky130_fd_sc_hd__o211a_1_1/X sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7385 sky130_fd_sc_hd__o221ai_1_0/a_295_297# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C7386 sky130_fd_sc_hd__dfrtn_1_16/a_805_47# sky130_fd_sc_hd__inv_1_25/A 0.00fF
C7387 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C7388 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C7389 sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C7390 sky130_fd_sc_hd__dfrtn_1_38/a_651_413# RESET_COUNTERn 0.01fF
C7391 sky130_fd_sc_hd__dfrtn_1_14/a_639_47# DOUT[18] 0.00fF
C7392 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__o211a_1_1/a_510_47# 0.00fF
C7393 CLK_REF sky130_fd_sc_hd__dfrtn_1_21/a_1217_47# 0.00fF
C7394 sky130_fd_sc_hd__dfrtn_1_14/a_651_413# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C7395 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# VDD 0.06fF
C7396 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C7397 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C7398 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C7399 sky130_fd_sc_hd__nand3b_1_1/Y sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C7400 sky130_fd_sc_hd__dfrtn_1_17/a_1462_47# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C7401 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__or2_2_0/B 0.02fF
C7402 sky130_fd_sc_hd__nor3_1_13/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7403 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C7404 sky130_fd_sc_hd__dfrtn_1_12/a_761_289# VDD 0.05fF
C7405 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_30/a_27_47# 0.00fF
C7406 sky130_fd_sc_hd__inv_1_28/A RESET_COUNTERn 0.15fF
C7407 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_10/a_805_47# 0.00fF
C7408 sky130_fd_sc_hd__dfrtn_1_39/a_651_413# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C7409 sky130_fd_sc_hd__dfrtn_1_17/a_543_47# sky130_fd_sc_hd__inv_1_28/Y 0.01fF
C7410 sky130_fd_sc_hd__inv_1_8/A DOUT[21] 0.23fF
C7411 sky130_fd_sc_hd__mux4_2_0/a_1064_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7412 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# DOUT[23] 0.00fF
C7413 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7414 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# DOUT[5] 0.00fF
C7415 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# -0.00fF
C7416 sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C7417 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_448_47# -0.00fF
C7418 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# DOUT[14] 0.00fF
C7419 sky130_fd_sc_hd__dfrtn_1_28/a_193_47# sky130_fd_sc_hd__inv_1_48/Y 0.06fF
C7420 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__o311a_1_0/a_585_47# 0.00fF
C7421 sky130_fd_sc_hd__dfrtn_1_18/a_651_413# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C7422 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C7423 sky130_fd_sc_hd__dfrtn_1_42/a_193_47# sky130_fd_sc_hd__nor3_2_2/A 0.53fF
C7424 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_2/a_639_47# 0.00fF
C7425 sky130_fd_sc_hd__dfrtn_1_26/a_639_47# RESET_COUNTERn 0.00fF
C7426 sky130_fd_sc_hd__nor3_1_20/a_193_297# DOUT[14] 0.00fF
C7427 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_34/a_761_289# 0.02fF
C7428 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C7429 sky130_fd_sc_hd__dfrtn_1_37/a_805_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C7430 sky130_fd_sc_hd__dfrtn_1_33/a_805_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C7431 DOUT[9] sky130_fd_sc_hd__nor3_1_2/a_109_297# 0.00fF
C7432 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__dfrtp_1_3/a_543_47# 0.01fF
C7433 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# sky130_fd_sc_hd__dfrtp_1_3/a_1283_21# 0.00fF
C7434 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_651_413# 0.00fF
C7435 sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C7436 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__dfrtp_1_3/a_448_47# 0.00fF
C7437 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C7438 sky130_fd_sc_hd__dfrtn_1_25/a_1217_47# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C7439 sky130_fd_sc_hd__dfrtn_1_16/a_1270_413# sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C7440 sky130_fd_sc_hd__dfrtn_1_11/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7441 sky130_fd_sc_hd__dfrtn_1_34/a_805_47# RESET_COUNTERn -0.00fF
C7442 sky130_fd_sc_hd__dfrtn_1_11/a_1462_47# VDD 0.00fF
C7443 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_21/a_761_289# 0.00fF
C7444 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_21/a_1270_413# 0.00fF
C7445 DOUT[13] sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C7446 sky130_fd_sc_hd__dfrtn_1_36/a_761_289# sky130_fd_sc_hd__inv_1_40/A 0.00fF
C7447 sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7448 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C7449 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__dfrtn_1_2/a_448_47# 0.00fF
C7450 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__dfrtn_1_37/a_27_47# 0.00fF
C7451 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__dfrtn_1_37/a_193_47# 0.01fF
C7452 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_37/a_543_47# 0.00fF
C7453 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_37/a_761_289# 0.01fF
C7454 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# sky130_fd_sc_hd__inv_1_48/A 0.01fF
C7455 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7456 DOUT[19] sky130_fd_sc_hd__nor3_2_3/B 0.11fF
C7457 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__nor3_2_0/A 0.01fF
C7458 sky130_fd_sc_hd__nor3_1_10/a_193_297# DOUT[19] 0.00fF
C7459 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C7460 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__dfrtn_1_2/a_543_47# 0.00fF
C7461 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_2/a_761_289# 0.00fF
C7462 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.01fF
C7463 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# 0.00fF
C7464 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# 0.01fF
C7465 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_35/a_651_413# 0.00fF
C7466 HEADER_2/a_508_138# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C7467 sky130_fd_sc_hd__dfrtn_1_34/a_1270_413# DONE 0.00fF
C7468 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__mux4_1_0/a_193_47# 0.00fF
C7469 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_24/a_193_47# -0.29fF
C7470 sky130_fd_sc_hd__o211a_1_1/a_510_47# DOUT[23] 0.00fF
C7471 sky130_fd_sc_hd__nor3_1_16/a_193_297# DOUT[4] 0.00fF
C7472 sky130_fd_sc_hd__nor3_1_12/a_193_297# DOUT[12] 0.00fF
C7473 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__inv_1_32/A 0.01fF
C7474 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C7475 DOUT[9] sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.00fF
C7476 sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C7477 sky130_fd_sc_hd__dfrtn_1_27/a_805_47# VDD 0.00fF
C7478 sky130_fd_sc_hd__dfrtn_1_27/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7479 sky130_fd_sc_hd__dfrtp_1_3/a_543_47# sky130_fd_sc_hd__or2_2_0/a_121_297# 0.00fF
C7480 sky130_fd_sc_hd__dfrtn_1_39/a_193_47# sky130_fd_sc_hd__inv_1_31/Y 0.01fF
C7481 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_18/a_805_47# 0.00fF
C7482 DOUT[1] sky130_fd_sc_hd__dfrtn_1_22/a_543_47# 0.00fF
C7483 sky130_fd_sc_hd__inv_1_47/Y SEL_CONV_TIME[2] 0.00fF
C7484 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# DOUT[21] 0.00fF
C7485 sky130_fd_sc_hd__dfrtn_1_21/a_193_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C7486 sky130_fd_sc_hd__nor3_2_3/a_281_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7487 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_805_47# -0.00fF
C7488 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__nor3_1_0/a_109_297# 0.00fF
C7489 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# DOUT[23] 0.00fF
C7490 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# DOUT[14] 0.00fF
C7491 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_3/a_27_47# 0.00fF
C7492 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_193_47# 0.00fF
C7493 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_761_289# 0.00fF
C7494 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__dfrtn_1_15/a_27_47# 0.00fF
C7495 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__inv_1_42/Y 0.27fF
C7496 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C7497 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C7498 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C7499 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C7500 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_12/A 0.00fF
C7501 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C7502 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__inv_1_49/A 0.05fF
C7503 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__nor3_1_0/a_193_297# 0.00fF
C7504 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7505 sky130_fd_sc_hd__dfrtn_1_36/a_761_289# VDD 0.05fF
C7506 sky130_fd_sc_hd__dfrtn_1_26/a_805_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C7507 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# 0.01fF
C7508 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_543_47# 0.00fF
C7509 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_761_289# 0.00fF
C7510 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# SEL_CONV_TIME[3] 0.00fF
C7511 sky130_fd_sc_hd__nor3_2_3/A RESET_COUNTERn 0.17fF
C7512 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7513 sky130_fd_sc_hd__dfrtn_1_26/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7514 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# VDD -0.00fF
C7515 sky130_fd_sc_hd__dfrtn_1_17/a_761_289# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C7516 sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C7517 sky130_fd_sc_hd__dfrtp_1_3/a_1462_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C7518 sky130_fd_sc_hd__inv_1_5/Y DOUT[14] 0.00fF
C7519 sky130_fd_sc_hd__dfrtn_1_34/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7520 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_27/a_448_47# 0.00fF
C7521 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# 0.00fF
C7522 sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__dfrtn_1_16/a_193_47# 0.00fF
C7523 sky130_fd_sc_hd__dfrtn_1_28/a_543_47# RESET_COUNTERn 0.01fF
C7524 sky130_fd_sc_hd__dfrtn_1_28/a_1270_413# DOUT[21] 0.00fF
C7525 sky130_fd_sc_hd__dfrtn_1_33/a_1462_47# DOUT[23] 0.00fF
C7526 sky130_fd_sc_hd__dfrtn_1_14/a_448_47# sky130_fd_sc_hd__nor3_1_1/a_193_297# 0.00fF
C7527 sky130_fd_sc_hd__dfrtn_1_14/a_651_413# sky130_fd_sc_hd__nor3_1_1/a_109_297# 0.00fF
C7528 sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C7529 sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C7530 sky130_fd_sc_hd__nor3_1_0/a_109_297# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C7531 sky130_fd_sc_hd__dfrtn_1_14/a_805_47# RESET_COUNTERn 0.00fF
C7532 sky130_fd_sc_hd__mux4_1_0/a_1478_413# SEL_CONV_TIME[0] 0.00fF
C7533 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_11/a_193_47# 0.00fF
C7534 DOUT[1] sky130_fd_sc_hd__nor3_2_2/a_27_297# 0.00fF
C7535 sky130_fd_sc_hd__dfrtn_1_42/a_1462_47# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C7536 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C7537 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C7538 sky130_fd_sc_hd__inv_1_25/A sky130_fd_sc_hd__nor3_2_3/B 0.08fF
C7539 sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C7540 sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C7541 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# SEL_CONV_TIME[2] 0.01fF
C7542 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# VIN 0.00fF
C7543 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C7544 sky130_fd_sc_hd__dfrtn_1_4/a_651_413# VIN 0.00fF
C7545 sky130_fd_sc_hd__dfrtn_1_14/a_639_47# DOUT[22] 0.00fF
C7546 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C7547 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C7548 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C7549 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C7550 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C7551 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C7552 sky130_fd_sc_hd__dfrtn_1_32/a_761_289# sky130_fd_sc_hd__inv_1_9/A 0.00fF
C7553 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__dfrtn_1_37/a_1462_47# 0.00fF
C7554 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# 0.00fF
C7555 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_37/a_639_47# 0.00fF
C7556 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# RESET_COUNTERn -0.01fF
C7557 DOUT[1] sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# 0.01fF
C7558 sky130_fd_sc_hd__dfrtn_1_18/a_761_289# DOUT[2] 0.01fF
C7559 sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7560 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__nor3_1_13/a_109_297# 0.00fF
C7561 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7562 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_25/a_651_413# 0.00fF
C7563 DOUT[2] sky130_fd_sc_hd__inv_1_40/Y 0.00fF
C7564 sky130_fd_sc_hd__dfrtn_1_22/a_1270_413# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C7565 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# -0.00fF
C7566 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7567 sky130_fd_sc_hd__inv_1_13/Y RESET_COUNTERn 0.03fF
C7568 sky130_fd_sc_hd__o221ai_1_0/a_213_123# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C7569 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C7570 sky130_fd_sc_hd__nor3_1_12/a_193_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7571 sky130_fd_sc_hd__or3b_2_0/a_388_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7572 sky130_fd_sc_hd__dfrtn_1_31/a_1108_47# SEL_CONV_TIME[1] 0.00fF
C7573 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_651_413# -0.00fF
C7574 sky130_fd_sc_hd__dfrtn_1_17/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_448_47# -0.00fF
C7575 sky130_fd_sc_hd__mux4_1_0/a_247_21# RESET_COUNTERn 0.03fF
C7576 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# RESET_COUNTERn 0.00fF
C7577 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_41/a_805_47# 0.00fF
C7578 sky130_fd_sc_hd__or3b_2_0/a_388_297# sky130_fd_sc_hd__dfrtn_1_31/a_193_47# 0.00fF
C7579 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_761_289# 0.00fF
C7580 sky130_fd_sc_hd__or3b_2_0/a_472_297# sky130_fd_sc_hd__dfrtn_1_31/a_27_47# 0.00fF
C7581 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_31/a_543_47# 0.00fF
C7582 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_19/a_651_413# 0.00fF
C7583 sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# DOUT[23] 0.00fF
C7584 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# DOUT[19] 0.00fF
C7585 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C7586 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__dfrtn_1_15/a_651_413# 0.00fF
C7587 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# 0.00fF
C7588 sky130_fd_sc_hd__dfrtn_1_25/a_1217_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C7589 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_639_47# 0.00fF
C7590 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C7591 sky130_fd_sc_hd__dfrtn_1_17/a_448_47# VDD 0.01fF
C7592 sky130_fd_sc_hd__dfrtn_1_28/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.05fF
C7593 SLC_0/a_264_22# outb 0.01fF
C7594 sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__inv_1_54/Y 0.00fF
C7595 sky130_fd_sc_hd__dfrtn_1_3/a_1270_413# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C7596 sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7597 sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7598 sky130_fd_sc_hd__inv_1_11/A sky130_fd_sc_hd__inv_1_12/A 0.00fF
C7599 sky130_fd_sc_hd__dfrtn_1_12/a_805_47# sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# 0.00fF
C7600 sky130_fd_sc_hd__dfrtn_1_32/a_27_47# sky130_fd_sc_hd__dfrtn_1_32/a_761_289# -0.00fF
C7601 sky130_fd_sc_hd__nor3_1_20/a_193_297# sky130_fd_sc_hd__dfrtn_1_22/a_1283_21# 0.00fF
C7602 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# 0.00fF
C7603 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_1462_47# 0.00fF
C7604 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__o2111a_2_0/a_566_47# 0.00fF
C7605 sky130_fd_sc_hd__nor3_2_3/a_281_297# sky130_fd_sc_hd__dfrtn_1_42/a_651_413# 0.00fF
C7606 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# 0.00fF
C7607 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C7608 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__inv_1_41/Y 0.01fF
C7609 sky130_fd_sc_hd__dfrtn_1_22/a_761_289# sky130_fd_sc_hd__inv_1_37/A 0.02fF
C7610 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C7611 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C7612 sky130_fd_sc_hd__nor3_1_7/a_193_297# DOUT[14] 0.00fF
C7613 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.01fF
C7614 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.01fF
C7615 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.01fF
C7616 sky130_fd_sc_hd__o211a_1_0/a_510_47# DOUT[15] 0.00fF
C7617 sky130_fd_sc_hd__o311a_1_0/a_266_47# SEL_CONV_TIME[0] 0.00fF
C7618 outb DOUT[10] 0.00fF
C7619 en VIN 1.38fF
C7620 sky130_fd_sc_hd__dfrtn_1_31/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7621 sky130_fd_sc_hd__conb_1_0/LO DOUT[23] 0.01fF
C7622 sky130_fd_sc_hd__dfrtn_1_31/a_1283_21# VDD 0.13fF
C7623 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_4/Y 0.01fF
C7624 sky130_fd_sc_hd__inv_1_38/Y sky130_fd_sc_hd__inv_1_40/A 0.00fF
C7625 sky130_fd_sc_hd__mux4_2_0/a_788_316# SEL_CONV_TIME[0] 0.02fF
C7626 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_11/a_1462_47# 0.00fF
C7627 sky130_fd_sc_hd__dfrtn_1_0/a_651_413# RESET_COUNTERn 0.00fF
C7628 sky130_fd_sc_hd__dfrtn_1_35/a_543_47# RESET_COUNTERn 0.01fF
C7629 sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C7630 sky130_fd_sc_hd__nor3_1_11/a_109_297# sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# 0.00fF
C7631 sky130_fd_sc_hd__nor3_1_11/a_193_297# sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# 0.00fF
C7632 sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C7633 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_543_47# -0.00fF
C7634 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# sky130_fd_sc_hd__dfrtn_1_31/a_761_289# -0.00fF
C7635 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C7636 sky130_fd_sc_hd__dfrtn_1_23/a_639_47# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C7637 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C7638 sky130_fd_sc_hd__or2b_1_0/a_301_297# SEL_CONV_TIME[1] 0.00fF
C7639 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# DOUT[3] 0.00fF
C7640 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_805_47# 0.00fF
C7641 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_30/a_651_413# 0.00fF
C7642 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# RESET_COUNTERn 0.00fF
C7643 sky130_fd_sc_hd__dfrtn_1_32/a_1462_47# sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# 0.00fF
C7644 sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# sky130_fd_sc_hd__dfrtn_1_36/a_1462_47# 0.00fF
C7645 sky130_fd_sc_hd__dfrtn_1_4/a_761_289# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C7646 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_19/a_448_47# 0.00fF
C7647 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__inv_1_31/A 0.00fF
C7648 sky130_fd_sc_hd__dfrtn_1_0/a_448_47# DOUT[22] 0.00fF
C7649 sky130_fd_sc_hd__dfrtn_1_20/a_1462_47# RESET_COUNTERn -0.00fF
C7650 sky130_fd_sc_hd__dfrtn_1_41/a_1270_413# SEL_CONV_TIME[0] 0.00fF
C7651 sky130_fd_sc_hd__dfrtn_1_21/a_761_289# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C7652 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__inv_1_43/Y 0.01fF
C7653 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C7654 sky130_fd_sc_hd__dfrtn_1_34/a_543_47# sky130_fd_sc_hd__o221ai_1_0/a_493_297# 0.00fF
C7655 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C7656 sky130_fd_sc_hd__dfrtp_1_2/a_805_47# sky130_fd_sc_hd__inv_1_29/Y 0.00fF
C7657 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__inv_1_2/A 0.01fF
C7658 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_18/a_543_47# 0.00fF
C7659 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_18/a_651_413# 0.00fF
C7660 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C7661 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_639_47# 0.00fF
C7662 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# 0.00fF
C7663 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_805_47# 0.00fF
C7664 sky130_fd_sc_hd__inv_1_30/A DOUT[2] 0.06fF
C7665 sky130_fd_sc_hd__dfrtn_1_42/a_651_413# sky130_fd_sc_hd__inv_1_25/A 0.00fF
C7666 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7667 sky130_fd_sc_hd__dfrtn_1_32/a_639_47# VDD 0.00fF
C7668 sky130_fd_sc_hd__dfrtn_1_32/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7669 sky130_fd_sc_hd__dfrtn_1_10/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7670 sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C7671 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# 0.00fF
C7672 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__inv_1_1/A 0.01fF
C7673 sky130_fd_sc_hd__dfrtn_1_3/a_651_413# DOUT[11] 0.00fF
C7674 sky130_fd_sc_hd__inv_1_33/A sky130_fd_sc_hd__inv_1_41/Y 0.07fF
C7675 sky130_fd_sc_hd__dfrtn_1_4/a_651_413# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C7676 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_1/a_761_289# -0.00fF
C7677 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# SEL_CONV_TIME[1] 0.03fF
C7678 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_38/a_805_47# 0.00fF
C7679 sky130_fd_sc_hd__dfrtn_1_36/a_651_413# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C7680 sky130_fd_sc_hd__inv_1_44/A RESET_COUNTERn 0.03fF
C7681 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C7682 sky130_fd_sc_hd__inv_1_6/Y DOUT[6] 0.04fF
C7683 sky130_fd_sc_hd__o311a_1_0/a_368_297# DOUT[21] 0.00fF
C7684 sky130_fd_sc_hd__or3_1_0/a_111_297# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C7685 sky130_fd_sc_hd__dfrtp_1_3/a_1108_47# sky130_fd_sc_hd__or2_2_0/A 0.01fF
C7686 sky130_fd_sc_hd__dfrtn_1_27/a_193_47# SEL_CONV_TIME[0] 0.00fF
C7687 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__inv_1_53/Y 0.01fF
C7688 sky130_fd_sc_hd__or2b_1_0/a_27_53# VDD 0.05fF
C7689 VDD sky130_fd_sc_hd__inv_1_38/Y 0.63fF
C7690 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# 0.00fF
C7691 sky130_fd_sc_hd__dfrtn_1_23/a_543_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C7692 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C7693 sky130_fd_sc_hd__inv_1_18/Y DOUT[12] 0.00fF
C7694 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_14/A 0.00fF
C7695 sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# sky130_fd_sc_hd__dfrtn_1_28/a_543_47# 0.00fF
C7696 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_36/a_761_289# 0.01fF
C7697 sky130_fd_sc_hd__nor3_1_15/a_109_297# DOUT[16] 0.00fF
C7698 sky130_fd_sc_hd__nor3_1_15/a_193_297# sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C7699 sky130_fd_sc_hd__dfrtn_1_34/a_639_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C7700 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C7701 sky130_fd_sc_hd__dfrtn_1_42/a_1108_47# sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C7702 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# sky130_fd_sc_hd__inv_1_14/A 0.10fF
C7703 sky130_fd_sc_hd__dfrtn_1_28/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7704 sky130_fd_sc_hd__dfrtn_1_4/a_543_47# DOUT[11] 0.00fF
C7705 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C7706 sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7707 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# DOUT[9] 0.00fF
C7708 sky130_fd_sc_hd__dfrtn_1_35/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7709 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# VDD 0.01fF
C7710 sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C7711 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__inv_1_33/A 0.02fF
C7712 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# RESET_COUNTERn 0.02fF
C7713 sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# 0.00fF
C7714 sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# 0.00fF
C7715 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_34/a_543_47# 0.00fF
C7716 sky130_fd_sc_hd__o311a_1_0/a_368_297# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C7717 DOUT[4] sky130_fd_sc_hd__dfrtn_1_30/a_651_413# 0.00fF
C7718 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__nor3_1_5/A 0.00fF
C7719 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__dfrtn_1_30/a_639_47# -0.00fF
C7720 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_805_47# 0.00fF
C7721 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C7722 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__dfrtn_1_5/a_448_47# 0.00fF
C7723 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C7724 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C7725 sky130_fd_sc_hd__o221ai_1_0/a_109_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C7726 sky130_fd_sc_hd__dfrtn_1_19/a_1283_21# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C7727 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfrtn_1_41/a_805_47# 0.00fF
C7728 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__inv_1_8/Y 0.01fF
C7729 sky130_fd_sc_hd__inv_1_14/A sky130_fd_sc_hd__inv_1_1/A 0.05fF
C7730 sky130_fd_sc_hd__dfrtn_1_3/a_805_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C7731 sky130_fd_sc_hd__dfrtn_1_38/a_805_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C7732 sky130_fd_sc_hd__dfrtn_1_28/a_805_47# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C7733 sky130_fd_sc_hd__dfrtn_1_25/a_651_413# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C7734 sky130_fd_sc_hd__dfrtn_1_32/a_543_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C7735 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__o211a_1_1/X 0.02fF
C7736 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# DOUT[21] 0.00fF
C7737 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_1/a_543_47# 0.00fF
C7738 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C7739 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C7740 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# DOUT[3] 0.00fF
C7741 sky130_fd_sc_hd__inv_1_37/A DOUT[15] 0.00fF
C7742 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_14/a_651_413# 0.00fF
C7743 sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# RESET_COUNTERn 0.00fF
C7744 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_25/a_543_47# 0.00fF
C7745 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_25/a_27_47# 0.00fF
C7746 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__dfrtn_1_25/a_193_47# 0.00fF
C7747 sky130_fd_sc_hd__dfrtp_1_3/a_639_47# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C7748 sky130_fd_sc_hd__dfrtp_1_3/a_805_47# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C7749 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_805_47# 0.00fF
C7750 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_639_47# 0.00fF
C7751 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C7752 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__mux4_2_0/a_193_369# 0.00fF
C7753 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__dfrtp_1_2/a_543_47# -0.00fF
C7754 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C7755 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C7756 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__inv_1_7/A 0.01fF
C7757 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7758 sky130_fd_sc_hd__dfrtn_1_4/a_448_47# sky130_fd_sc_hd__inv_1_7/A 0.01fF
C7759 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# CLK_REF 0.00fF
C7760 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__nor3_1_19/Y 0.01fF
C7761 sky130_fd_sc_hd__dfrtp_1_3/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7762 sky130_fd_sc_hd__dfrtp_1_3/a_639_47# VDD 0.00fF
C7763 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.01fF
C7764 sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# SEL_CONV_TIME[1] 0.00fF
C7765 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# VDD 0.19fF
C7766 sky130_fd_sc_hd__dfrtn_1_21/a_805_47# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C7767 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C7768 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C7769 sky130_fd_sc_hd__dfrtn_1_28/a_761_289# sky130_fd_sc_hd__inv_1_48/A 0.02fF
C7770 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C7771 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__dfrtn_1_24/a_193_47# 0.00fF
C7772 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__dfrtn_1_24/a_761_289# 0.00fF
C7773 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# 0.00fF
C7774 sky130_fd_sc_hd__dfrtn_1_27/a_1462_47# SEL_CONV_TIME[0] 0.00fF
C7775 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C7776 DOUT[4] sky130_fd_sc_hd__dfrtn_1_34/a_543_47# 0.01fF
C7777 sky130_fd_sc_hd__dfrtn_1_25/a_1462_47# sky130_fd_sc_hd__dfrtn_1_28/a_448_47# 0.00fF
C7778 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__dfrtp_1_1/D 0.00fF
C7779 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__o211a_1_1/a_510_47# 0.00fF
C7780 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C7781 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# sky130_fd_sc_hd__inv_1_40/A 0.01fF
C7782 sky130_fd_sc_hd__inv_1_32/A RESET_COUNTERn 0.30fF
C7783 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_448_47# -0.00fF
C7784 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_651_413# -0.00fF
C7785 sky130_fd_sc_hd__inv_1_44/A SEL_CONV_TIME[3] 0.01fF
C7786 sky130_fd_sc_hd__inv_1_44/Y DOUT[21] 0.03fF
C7787 sky130_fd_sc_hd__dfrtn_1_11/a_1270_413# RESET_COUNTERn 0.00fF
C7788 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# DOUT[23] 0.00fF
C7789 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_10/a_543_47# 0.00fF
C7790 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# DOUT[19] 0.00fF
C7791 sky130_fd_sc_hd__dfrtn_1_35/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7792 sky130_fd_sc_hd__dfrtn_1_8/a_543_47# DOUT[12] 0.00fF
C7793 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__nor3_2_0/A 0.54fF
C7794 sky130_fd_sc_hd__nor3_2_0/a_281_297# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C7795 sky130_fd_sc_hd__inv_1_19/A sky130_fd_sc_hd__inv_1_23/A 0.13fF
C7796 sky130_fd_sc_hd__nor3_1_0/a_109_297# DOUT[17] 0.00fF
C7797 sky130_fd_sc_hd__nor3_1_11/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7798 sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7799 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__inv_1_53/A 0.01fF
C7800 sky130_fd_sc_hd__dfrtn_1_29/a_805_47# VDD 0.00fF
C7801 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__dfrtp_1_3/a_761_289# -0.00fF
C7802 sky130_fd_sc_hd__inv_1_13/Y DOUT[10] 0.01fF
C7803 sky130_fd_sc_hd__dfrtp_1_1/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7804 CLK_REF sky130_fd_sc_hd__dfrtn_1_19/a_543_47# 0.01fF
C7805 sky130_fd_sc_hd__nand2_1_2/a_113_47# SEL_CONV_TIME[0] 0.00fF
C7806 sky130_fd_sc_hd__dfrtp_1_2/a_805_47# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.00fF
C7807 sky130_fd_sc_hd__nor3_1_3/a_109_297# VDD 0.00fF
C7808 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C7809 sky130_fd_sc_hd__dfrtn_1_18/a_761_289# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C7810 sky130_fd_sc_hd__dfrtn_1_20/a_1270_413# sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.00fF
C7811 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__dfrtn_1_29/a_761_289# 0.00fF
C7812 sky130_fd_sc_hd__nor3_1_16/a_109_297# sky130_fd_sc_hd__dfrtn_1_35/a_1283_21# 0.00fF
C7813 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# DOUT[2] 0.01fF
C7814 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__nor3_2_1/A 0.12fF
C7815 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C7816 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_34/a_543_47# 0.00fF
C7817 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__o211a_1_0/a_215_47# 0.00fF
C7818 sky130_fd_sc_hd__dfrtn_1_23/a_1270_413# sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C7819 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# 0.00fF
C7820 sky130_fd_sc_hd__dfrtn_1_23/a_543_47# sky130_fd_sc_hd__dfrtn_1_36/a_448_47# 0.00fF
C7821 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__o211a_1_0/a_297_297# 0.00fF
C7822 sky130_fd_sc_hd__dfrtn_1_23/a_639_47# sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C7823 sky130_fd_sc_hd__inv_1_41/Y sky130_fd_sc_hd__o2111a_2_0/X 0.03fF
C7824 SEL_CONV_TIME[2] sky130_fd_sc_hd__inv_1_44/A 0.00fF
C7825 sky130_fd_sc_hd__o311a_1_0/A3 sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C7826 SEL_CONV_TIME[1] sky130_fd_sc_hd__inv_1_48/Y 0.01fF
C7827 sky130_fd_sc_hd__dfrtn_1_27/a_448_47# RESET_COUNTERn 0.01fF
C7828 sky130_fd_sc_hd__inv_1_43/Y sky130_fd_sc_hd__inv_1_43/A 0.09fF
C7829 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C7830 sky130_fd_sc_hd__dfrtn_1_27/a_1217_47# DOUT[21] 0.00fF
C7831 sky130_fd_sc_hd__dfrtn_1_38/a_651_413# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C7832 sky130_fd_sc_hd__dfrtn_1_35/a_651_413# sky130_fd_sc_hd__inv_1_38/A 0.00fF
C7833 sky130_fd_sc_hd__nor3_1_18/a_193_297# RESET_COUNTERn 0.00fF
C7834 sky130_fd_sc_hd__dfrtn_1_11/a_805_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C7835 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__inv_1_41/Y -0.01fF
C7836 sky130_fd_sc_hd__dfrtn_1_9/a_761_289# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C7837 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# VDD 0.09fF
C7838 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__dfrtn_1_25/a_639_47# 0.00fF
C7839 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_35/a_27_47# 0.00fF
C7840 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_32/a_639_47# 0.00fF
C7841 sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C7842 sky130_fd_sc_hd__nor3_2_0/a_281_297# sky130_fd_sc_hd__dfrtn_1_12/a_543_47# 0.00fF
C7843 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__dfrtn_1_34/a_761_289# -0.00fF
C7844 VDD DOUT[18] 1.29fF
C7845 DOUT[13] sky130_fd_sc_hd__dfrtn_1_30/a_761_289# 0.01fF
C7846 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# sky130_fd_sc_hd__mux4_2_0/a_872_316# 0.00fF
C7847 sky130_fd_sc_hd__dfrtn_1_37/a_1462_47# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C7848 sky130_fd_sc_hd__dfrtn_1_37/a_1270_413# sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C7849 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# sky130_fd_sc_hd__mux4_2_0/a_1060_369# 0.00fF
C7850 sky130_fd_sc_hd__dfrtn_1_37/a_805_47# sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.00fF
C7851 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# sky130_fd_sc_hd__mux4_2_0/a_193_47# 0.00fF
C7852 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C7853 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# sky130_fd_sc_hd__mux4_2_0/a_600_345# 0.00fF
C7854 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C7855 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_761_289# 0.00fF
C7856 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# sky130_fd_sc_hd__mux4_2_0/a_397_47# 0.00fF
C7857 sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# DOUT[2] 0.00fF
C7858 sky130_fd_sc_hd__mux4_2_0/a_872_316# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7859 sky130_fd_sc_hd__dfrtn_1_10/a_805_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C7860 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# sky130_fd_sc_hd__inv_1_32/A 0.03fF
C7861 sky130_fd_sc_hd__dfrtn_1_36/a_543_47# DOUT[21] 0.01fF
C7862 sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C7863 sky130_fd_sc_hd__inv_1_45/Y DOUT[23] 0.00fF
C7864 sky130_fd_sc_hd__nand3b_1_1/Y sky130_fd_sc_hd__nor3_1_19/Y 0.45fF
C7865 sky130_fd_sc_hd__dfrtn_1_21/a_761_289# VDD 0.05fF
C7866 sky130_fd_sc_hd__nor3_2_3/a_281_297# DOUT[2] 0.00fF
C7867 sky130_fd_sc_hd__o221ai_1_0/a_493_297# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C7868 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__or2_2_0/B 0.03fF
C7869 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# RESET_COUNTERn 0.00fF
C7870 sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C7871 sky130_fd_sc_hd__dfrtn_1_33/a_651_413# sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# 0.00fF
C7872 sky130_fd_sc_hd__dfrtn_1_33/a_448_47# sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# 0.00fF
C7873 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# 0.00fF
C7874 sky130_fd_sc_hd__dfrtn_1_14/a_543_47# sky130_fd_sc_hd__inv_1_0/Y 0.01fF
C7875 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C7876 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C7877 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# sky130_fd_sc_hd__nor3_1_1/a_193_297# 0.00fF
C7878 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# VDD 0.04fF
C7879 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__inv_1_38/Y 0.12fF
C7880 sky130_fd_sc_hd__dfrtn_1_34/a_1462_47# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C7881 sky130_fd_sc_hd__dfrtn_1_22/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7882 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__nor3_1_1/a_109_297# 0.00fF
C7883 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_651_413# -0.00fF
C7884 sky130_fd_sc_hd__dfrtn_1_38/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_448_47# -0.00fF
C7885 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_21/a_1462_47# 0.00fF
C7886 sky130_fd_sc_hd__dfrtn_1_22/a_1217_47# VDD 0.00fF
C7887 DOUT[1] sky130_fd_sc_hd__dfrtn_1_42/a_639_47# 0.00fF
C7888 sky130_fd_sc_hd__nor3_1_12/a_109_297# sky130_fd_sc_hd__dfrtn_1_8/a_543_47# 0.00fF
C7889 sky130_fd_sc_hd__nor3_1_12/a_193_297# sky130_fd_sc_hd__dfrtn_1_8/a_761_289# 0.00fF
C7890 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7891 sky130_fd_sc_hd__dfrtn_1_12/a_639_47# RESET_COUNTERn 0.00fF
C7892 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__inv_1_1/A 0.02fF
C7893 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__dfrtn_1_25/a_543_47# 0.00fF
C7894 sky130_fd_sc_hd__nand3b_1_0/a_316_47# sky130_fd_sc_hd__dfrtn_1_25/a_193_47# 0.00fF
C7895 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__inv_1_53/Y 0.04fF
C7896 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# 0.00fF
C7897 sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# sky130_fd_sc_hd__inv_1_53/Y 0.01fF
C7898 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__or2b_1_0/X 0.01fF
C7899 sky130_fd_sc_hd__dfrtn_1_23/a_1462_47# sky130_fd_sc_hd__inv_1_40/A 0.00fF
C7900 sky130_fd_sc_hd__dfrtp_1_0/a_761_289# sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# 0.00fF
C7901 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# 0.00fF
C7902 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# sky130_fd_sc_hd__dfrtp_1_1/a_193_47# 0.00fF
C7903 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__dfrtp_1_1/a_651_413# 0.00fF
C7904 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__mux4_2_0/a_872_316# 0.00fF
C7905 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__mux4_2_0/a_600_345# 0.00fF
C7906 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# 0.00fF
C7907 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__nor3_1_4/A 0.02fF
C7908 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_1270_413# 0.00fF
C7909 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C7910 sky130_fd_sc_hd__nor2_1_0/a_109_297# SEL_CONV_TIME[0] 0.00fF
C7911 sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C7912 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C7913 sky130_fd_sc_hd__mux4_2_0/a_1279_413# SEL_CONV_TIME[3] 0.00fF
C7914 sky130_fd_sc_hd__dfrtn_1_16/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7915 sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.03fF
C7916 sky130_fd_sc_hd__dfrtn_1_16/a_639_47# VDD 0.00fF
C7917 sky130_fd_sc_hd__dfrtn_1_8/a_1108_47# VDD 0.07fF
C7918 sky130_fd_sc_hd__dfrtn_1_8/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C7919 sky130_fd_sc_hd__dfrtn_1_3/a_1270_413# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C7920 sky130_fd_sc_hd__nor3_1_19/Y sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C7921 sky130_fd_sc_hd__nor3_2_2/A sky130_fd_sc_hd__nor3_2_3/A 0.02fF
C7922 sky130_fd_sc_hd__inv_1_25/A DOUT[2] 0.19fF
C7923 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__inv_1_49/A 0.04fF
C7924 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# -0.00fF
C7925 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__dfrtn_1_29/a_543_47# -0.00fF
C7926 sky130_fd_sc_hd__inv_1_32/A SEL_CONV_TIME[3] 0.01fF
C7927 sky130_fd_sc_hd__dfrtn_1_7/a_448_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C7928 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__inv_1_7/A 0.45fF
C7929 sky130_fd_sc_hd__a221oi_4_0/a_471_297# RESET_COUNTERn 0.00fF
C7930 sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C7931 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_20/a_651_413# 0.00fF
C7932 sky130_fd_sc_hd__dfrtp_1_2/a_805_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C7933 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__inv_1_30/Y 0.05fF
C7934 sky130_fd_sc_hd__dfrtn_1_31/a_448_47# SEL_CONV_TIME[0] 0.00fF
C7935 sky130_fd_sc_hd__dfrtp_1_0/a_1217_47# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C7936 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C7937 sky130_fd_sc_hd__inv_1_3/A DOUT[8] 0.01fF
C7938 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C7939 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C7940 sky130_fd_sc_hd__or3b_2_0/a_176_21# RESET_COUNTERn 0.04fF
C7941 sky130_fd_sc_hd__inv_1_33/A sky130_fd_sc_hd__inv_1_53/Y 0.01fF
C7942 DOUT[23] sky130_fd_sc_hd__or3_1_0/C 0.00fF
C7943 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7944 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__or3_1_0/C 0.03fF
C7945 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.00fF
C7946 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# 0.00fF
C7947 sky130_fd_sc_hd__dfrtn_1_23/a_1462_47# VDD 0.00fF
C7948 sky130_fd_sc_hd__dfrtn_1_12/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C7949 DONE SEL_CONV_TIME[1] 0.05fF
C7950 sky130_fd_sc_hd__inv_1_32/A SEL_CONV_TIME[2] 0.29fF
C7951 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__mux4_2_0/a_193_369# 0.00fF
C7952 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_1462_47# 0.00fF
C7953 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_38/a_651_413# 0.00fF
C7954 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# 0.00fF
C7955 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# 0.00fF
C7956 sky130_fd_sc_hd__dfrtn_1_7/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7957 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__or3b_2_0/a_388_297# 0.00fF
C7958 sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# VDD 0.00fF
C7959 sky130_fd_sc_hd__dfrtn_1_17/a_761_289# RESET_COUNTERn 0.02fF
C7960 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# DOUT[14] 0.01fF
C7961 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C7962 sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C7963 sky130_fd_sc_hd__dfrtn_1_36/a_639_47# RESET_COUNTERn 0.00fF
C7964 sky130_fd_sc_hd__dfrtn_1_3/a_651_413# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C7965 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C7966 sky130_fd_sc_hd__dfrtp_1_0/a_1217_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C7967 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_7/A 0.02fF
C7968 DOUT[9] sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C7969 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C7970 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__inv_1_0/Y 0.01fF
C7971 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__inv_1_11/Y 0.14fF
C7972 sky130_fd_sc_hd__nor3_2_3/C DOUT[8] 0.05fF
C7973 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_543_47# 0.00fF
C7974 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C7975 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_761_289# 0.00fF
C7976 sky130_fd_sc_hd__mux4_2_0/a_872_316# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C7977 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__or2_2_0/A 0.00fF
C7978 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C7979 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C7980 sky130_fd_sc_hd__dfrtn_1_18/a_448_47# sky130_fd_sc_hd__inv_1_35/A 0.00fF
C7981 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# RESET_COUNTERn 0.05fF
C7982 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C7983 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__inv_1_13/Y 0.01fF
C7984 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__nor3_1_4/A 0.22fF
C7985 sky130_fd_sc_hd__or2_2_0/a_39_297# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C7986 sky130_fd_sc_hd__dfrtn_1_27/a_639_47# DOUT[23] 0.00fF
C7987 DOUT[4] sky130_fd_sc_hd__inv_1_47/A 0.01fF
C7988 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# 0.00fF
C7989 sky130_fd_sc_hd__nor3_1_13/a_193_297# sky130_fd_sc_hd__dfrtn_1_10/a_193_47# 0.00fF
C7990 VDD DOUT[22] 2.22fF
C7991 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C7992 sky130_fd_sc_hd__dfrtp_1_1/a_639_47# DOUT[0] 0.00fF
C7993 sky130_fd_sc_hd__dfrtn_1_4/a_543_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C7994 CLK_REF sky130_fd_sc_hd__o211a_1_1/a_510_47# 0.00fF
C7995 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C7996 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C7997 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# SEL_CONV_TIME[1] 0.01fF
C7998 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_805_47# 0.00fF
C7999 sky130_fd_sc_hd__dfrtn_1_25/a_805_47# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C8000 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# sky130_fd_sc_hd__dfrtn_1_27/a_1270_413# 0.00fF
C8001 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_639_47# 0.00fF
C8002 sky130_fd_sc_hd__dfrtn_1_25/a_639_47# sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.00fF
C8003 sky130_fd_sc_hd__inv_1_14/A sky130_fd_sc_hd__nor3_2_0/A 0.39fF
C8004 sky130_fd_sc_hd__dfrtn_1_33/a_1108_47# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C8005 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C8006 SEL_CONV_TIME[1] sky130_fd_sc_hd__nor3_2_3/B 0.10fF
C8007 sky130_fd_sc_hd__o311a_1_0/a_81_21# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C8008 sky130_fd_sc_hd__nor3_1_4/a_193_297# DOUT[8] 0.00fF
C8009 sky130_fd_sc_hd__nor3_1_4/a_109_297# RESET_COUNTERn 0.00fF
C8010 sky130_fd_sc_hd__dfrtn_1_42/a_1270_413# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C8011 sky130_fd_sc_hd__inv_1_14/A DOUT[17] 0.00fF
C8012 sky130_fd_sc_hd__mux4_2_0/a_193_369# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C8013 DOUT[9] sky130_fd_sc_hd__inv_1_15/A 0.01fF
C8014 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_14/a_193_47# 0.00fF
C8015 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C8016 sky130_fd_sc_hd__dfrtn_1_34/a_1217_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C8017 sky130_fd_sc_hd__or3_1_0/X sky130_fd_sc_hd__inv_1_44/A 0.02fF
C8018 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C8019 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C8020 sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# RESET_COUNTERn 0.01fF
C8021 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# SEL_CONV_TIME[0] 0.02fF
C8022 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_33/a_193_47# 0.00fF
C8023 sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__dfrtn_1_33/a_27_47# 0.00fF
C8024 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C8025 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__dfrtn_1_34/a_651_413# 0.00fF
C8026 sky130_fd_sc_hd__nor3_2_1/a_27_297# RESET_COUNTERn 0.00fF
C8027 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__dfrtn_1_14/a_761_289# -0.00fF
C8028 sky130_fd_sc_hd__dfrtn_1_8/a_1283_21# sky130_fd_sc_hd__inv_1_9/Y 0.00fF
C8029 sky130_fd_sc_hd__dfrtn_1_28/a_543_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C8030 sky130_fd_sc_hd__dfrtp_1_2/a_639_47# CLK_REF 0.00fF
C8031 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C8032 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8033 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__dfrtn_1_22/a_448_47# -0.00fF
C8034 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# sky130_fd_sc_hd__dfrtn_1_22/a_1108_47# -0.00fF
C8035 sky130_fd_sc_hd__nor3_1_14/a_109_297# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C8036 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__or3b_2_0/a_472_297# 0.00fF
C8037 sky130_fd_sc_hd__mux4_1_0/a_27_413# DOUT[2] 0.00fF
C8038 sky130_fd_sc_hd__dfrtn_1_36/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8039 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# 0.00fF
C8040 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_23/a_193_47# 0.00fF
C8041 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C8042 sky130_fd_sc_hd__nand3b_1_1/a_53_93# SEL_CONV_TIME[1] 0.08fF
C8043 sky130_fd_sc_hd__dfrtn_1_24/a_1270_413# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C8044 sky130_fd_sc_hd__or3_1_0/a_29_53# SEL_CONV_TIME[1] 0.02fF
C8045 sky130_fd_sc_hd__a221oi_4_0/a_471_297# SEL_CONV_TIME[3] 0.02fF
C8046 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__inv_1_47/A 0.02fF
C8047 sky130_fd_sc_hd__or2b_1_0/a_301_297# DOUT[21] 0.00fF
C8048 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_1/A 0.00fF
C8049 sky130_fd_sc_hd__dfrtn_1_7/a_805_47# DOUT[14] 0.00fF
C8050 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# VDD 0.09fF
C8051 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_43/Y 0.01fF
C8052 DOUT[23] sky130_fd_sc_hd__or2_2_0/A 0.00fF
C8053 DOUT[1] sky130_fd_sc_hd__inv_1_39/Y 0.14fF
C8054 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C8055 sky130_fd_sc_hd__inv_1_52/Y DOUT[21] 0.01fF
C8056 sky130_fd_sc_hd__dfrtn_1_25/a_1462_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C8057 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# 0.00fF
C8058 sky130_fd_sc_hd__nor3_1_10/a_109_297# VDD 0.00fF
C8059 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C8060 sky130_fd_sc_hd__dfrtn_1_39/a_1270_413# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C8061 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# VDD 0.05fF
C8062 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# sky130_fd_sc_hd__inv_1_1/A 0.16fF
C8063 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__mux4_2_0/a_1281_47# 0.00fF
C8064 sky130_fd_sc_hd__inv_1_27/A SEL_CONV_TIME[0] 0.09fF
C8065 sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C8066 sky130_fd_sc_hd__nor3_1_3/a_109_297# DOUT[3] 0.00fF
C8067 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# RESET_COUNTERn 0.01fF
C8068 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C8069 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.01fF
C8070 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C8071 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C8072 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_1462_47# 0.00fF
C8073 sky130_fd_sc_hd__inv_1_19/A DOUT[10] 0.01fF
C8074 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C8075 sky130_fd_sc_hd__inv_1_13/Y sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C8076 sky130_fd_sc_hd__dfrtn_1_19/a_1108_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C8077 sky130_fd_sc_hd__dfrtn_1_0/a_1217_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C8078 DOUT[4] sky130_fd_sc_hd__dfrtn_1_35/a_651_413# 0.00fF
C8079 sky130_fd_sc_hd__dfrtn_1_11/a_1462_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C8080 sky130_fd_sc_hd__nor3_1_3/a_109_297# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C8081 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# DOUT[21] 0.01fF
C8082 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# 0.00fF
C8083 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# 0.00fF
C8084 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# 0.00fF
C8085 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# 0.00fF
C8086 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_31/a_543_47# 0.00fF
C8087 sky130_fd_sc_hd__a221oi_4_0/a_471_297# SEL_CONV_TIME[2] 0.00fF
C8088 sky130_fd_sc_hd__or2b_1_0/a_301_297# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C8089 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C8090 sky130_fd_sc_hd__dfrtn_1_31/a_1217_47# RESET_COUNTERn 0.00fF
C8091 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_37/a_27_47# 0.00fF
C8092 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C8093 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.00fF
C8094 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__dfrtn_1_26/a_761_289# 0.00fF
C8095 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__dfrtn_1_26/a_543_47# 0.00fF
C8096 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# 0.00fF
C8097 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__dfrtn_1_28/a_193_47# 0.00fF
C8098 sky130_fd_sc_hd__inv_1_9/Y RESET_COUNTERn 0.22fF
C8099 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_12/a_448_47# 0.00fF
C8100 sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C8101 sky130_fd_sc_hd__dfrtn_1_32/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8102 sky130_fd_sc_hd__dfrtn_1_25/a_448_47# SEL_CONV_TIME[1] 0.00fF
C8103 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__nor3_1_5/A 0.28fF
C8104 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C8105 sky130_fd_sc_hd__dfrtn_1_11/a_639_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C8106 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C8107 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# 0.00fF
C8108 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_8/a_1108_47# 0.01fF
C8109 sky130_fd_sc_hd__dfrtn_1_19/a_761_289# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C8110 sky130_fd_sc_hd__dfrtn_1_20/a_805_47# DOUT[2] 0.00fF
C8111 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# sky130_fd_sc_hd__dfrtn_1_16/a_761_289# -0.00fF
C8112 sky130_fd_sc_hd__nor3_1_9/a_109_297# VDD 0.00fF
C8113 DOUT[5] DOUT[18] 0.03fF
C8114 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__dfrtn_1_23/a_651_413# 0.00fF
C8115 sky130_fd_sc_hd__dfrtn_1_22/a_651_413# sky130_fd_sc_hd__dfrtn_1_23/a_27_47# 0.00fF
C8116 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# sky130_fd_sc_hd__dfrtn_1_23/a_448_47# 0.00fF
C8117 sky130_fd_sc_hd__dfrtn_1_22/a_448_47# sky130_fd_sc_hd__dfrtn_1_23/a_193_47# 0.00fF
C8118 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# DOUT[3] 0.00fF
C8119 sky130_fd_sc_hd__inv_1_53/A sky130_fd_sc_hd__inv_1_44/A 0.00fF
C8120 sky130_fd_sc_hd__dfrtn_1_31/a_639_47# DONE 0.00fF
C8121 sky130_fd_sc_hd__o221ai_1_0/a_109_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C8122 sky130_fd_sc_hd__mux4_2_0/a_1281_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C8123 sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C8124 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__o311a_1_0/A3 0.03fF
C8125 sky130_fd_sc_hd__dfrtn_1_38/a_448_47# sky130_fd_sc_hd__inv_1_27/Y 0.00fF
C8126 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# 0.00fF
C8127 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__dfrtn_1_16/a_193_47# 0.00fF
C8128 sky130_fd_sc_hd__nor3_2_2/a_281_297# sky130_fd_sc_hd__dfrtn_1_16/a_27_47# 0.00fF
C8129 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__inv_1_2/A 0.02fF
C8130 sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# SEL_CONV_TIME[0] 0.00fF
C8131 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_33/a_639_47# 0.00fF
C8132 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__dfrtn_1_33/a_543_47# 0.00fF
C8133 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__dfrtn_1_33/a_1270_413# 0.00fF
C8134 sky130_fd_sc_hd__nand2_1_1/Y SEL_CONV_TIME[1] 0.00fF
C8135 sky130_fd_sc_hd__nand3b_1_1/Y SEL_CONV_TIME[0] 0.04fF
C8136 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C8137 VDD sky130_fd_sc_hd__inv_1_6/A 0.77fF
C8138 sky130_fd_sc_hd__dfrtp_1_3/a_1108_47# RESET_COUNTERn 0.02fF
C8139 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1_6/a_193_47# -0.14fF
C8140 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__o211a_1_1/a_510_47# 0.00fF
C8141 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__o211a_1_1/a_297_297# 0.00fF
C8142 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__o211a_1_1/a_215_47# 0.00fF
C8143 sky130_fd_sc_hd__nor3_1_4/a_109_297# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C8144 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C8145 sky130_fd_sc_hd__or3_1_0/a_111_297# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C8146 sky130_fd_sc_hd__dfrtn_1_10/a_805_47# outb 0.00fF
C8147 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.01fF
C8148 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_23/a_1462_47# 0.00fF
C8149 sky130_fd_sc_hd__dfrtp_1_1/a_448_47# sky130_fd_sc_hd__o211a_1_1/X 0.00fF
C8150 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8151 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8152 sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# VDD 0.07fF
C8153 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C8154 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__dfrtn_1_3/a_27_47# 0.01fF
C8155 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__dfrtn_1_3/a_761_289# 0.00fF
C8156 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_3/a_193_47# 0.00fF
C8157 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_3/a_543_47# 0.00fF
C8158 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C8159 sky130_fd_sc_hd__dfrtn_1_12/a_1217_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C8160 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__inv_1_46/Y 0.00fF
C8161 sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# sky130_fd_sc_hd__inv_1_35/Y 0.00fF
C8162 sky130_fd_sc_hd__dfrtn_1_3/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8163 CLK_REF sky130_fd_sc_hd__conb_1_0/LO 0.00fF
C8164 sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C8165 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C8166 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# DOUT[2] 0.01fF
C8167 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# 0.00fF
C8168 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__dfrtp_1_2/a_543_47# 0.00fF
C8169 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__dfrtp_1_2/a_651_413# 0.00fF
C8170 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C8171 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C8172 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C8173 DOUT[1] sky130_fd_sc_hd__nor3_2_3/a_27_297# 0.00fF
C8174 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C8175 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# 0.00fF
C8176 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_805_47# 0.00fF
C8177 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C8178 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# 0.00fF
C8179 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# sky130_fd_sc_hd__inv_1_44/Y 0.01fF
C8180 sky130_fd_sc_hd__nor3_1_15/a_109_297# RESET_COUNTERn 0.00fF
C8181 sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C8182 sky130_fd_sc_hd__nor3_1_7/a_109_297# DOUT[9] 0.00fF
C8183 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C8184 sky130_fd_sc_hd__dfrtn_1_42/a_448_47# VDD 0.04fF
C8185 sky130_fd_sc_hd__inv_1_45/A DOUT[23] 0.00fF
C8186 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# DOUT[14] 0.00fF
C8187 sky130_fd_sc_hd__o311a_1_0/a_81_21# sky130_fd_sc_hd__o2111a_2_0/X 0.01fF
C8188 SEL_CONV_TIME[0] sky130_fd_sc_hd__inv_1_51/Y 0.01fF
C8189 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C8190 sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# DOUT[21] 0.00fF
C8191 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# RESET_COUNTERn 0.00fF
C8192 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C8193 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_44/A 0.00fF
C8194 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_25/a_193_47# 0.00fF
C8195 sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C8196 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_36/a_448_47# 0.00fF
C8197 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_761_289# 0.00fF
C8198 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C8199 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C8200 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.01fF
C8201 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C8202 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# VDD 0.00fF
C8203 sky130_fd_sc_hd__nor3_1_3/a_109_297# DOUT[20] 0.00fF
C8204 sky130_fd_sc_hd__dfrtn_1_4/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8205 sky130_fd_sc_hd__dfrtn_1_9/a_805_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C8206 sky130_fd_sc_hd__dfrtn_1_4/a_805_47# VDD 0.00fF
C8207 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_1/a_27_47# 0.01fF
C8208 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# 0.00fF
C8209 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# 0.00fF
C8210 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__mux4_2_0/a_193_369# 0.00fF
C8211 HEADER_1/a_508_138# RESET_COUNTERn 0.00fF
C8212 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C8213 sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# DOUT[3] 0.00fF
C8214 sky130_fd_sc_hd__dfrtn_1_19/a_193_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C8215 sky130_fd_sc_hd__inv_1_54/Y SEL_CONV_TIME[0] 0.00fF
C8216 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__or2_2_0/a_121_297# 0.00fF
C8217 SLC_0/a_438_293# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8218 SLC_0/a_919_243# VDD 0.10fF
C8219 sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C8220 sky130_fd_sc_hd__dfrtp_1_3/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8221 sky130_fd_sc_hd__dfrtn_1_16/a_761_289# DOUT[15] 0.01fF
C8222 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# sky130_fd_sc_hd__inv_1_43/A 0.01fF
C8223 sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C8224 sky130_fd_sc_hd__dfrtn_1_23/a_761_289# DOUT[21] 0.00fF
C8225 sky130_fd_sc_hd__dfrtn_1_8/a_27_47# sky130_fd_sc_hd__dfrtn_1_8/a_1108_47# -0.00fF
C8226 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C8227 sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C8228 sky130_fd_sc_hd__nand3b_1_0/a_316_47# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C8229 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__dfrtn_1_21/a_543_47# -0.00fF
C8230 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__dfrtn_1_7/a_193_47# 0.00fF
C8231 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# 0.00fF
C8232 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__dfrtn_1_7/a_543_47# 0.00fF
C8233 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C8234 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_3/a_1270_413# 0.00fF
C8235 DOUT[4] sky130_fd_sc_hd__dfrtn_1_12/a_761_289# 0.00fF
C8236 sky130_fd_sc_hd__dfrtn_1_12/a_761_289# sky130_fd_sc_hd__inv_1_0/Y 0.02fF
C8237 sky130_fd_sc_hd__nor3_2_2/a_281_297# DOUT[15] 0.02fF
C8238 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_0/a_639_47# 0.00fF
C8239 sky130_fd_sc_hd__mux4_2_0/a_1279_413# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C8240 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__dfrtn_1_28/a_805_47# -0.00fF
C8241 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8242 sky130_fd_sc_hd__dfrtp_1_0/a_1270_413# VDD 0.00fF
C8243 sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C8244 VDD out 3.63fF
C8245 sky130_fd_sc_hd__inv_1_54/A VDD 0.51fF
C8246 sky130_fd_sc_hd__inv_1_50/Y sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8247 sky130_fd_sc_hd__inv_1_32/A sky130_fd_sc_hd__inv_1_53/A 0.03fF
C8248 sky130_fd_sc_hd__inv_1_36/Y sky130_fd_sc_hd__inv_1_9/A 0.02fF
C8249 VDD sky130_fd_sc_hd__inv_1_48/A 0.92fF
C8250 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C8251 sky130_fd_sc_hd__inv_1_4/A DOUT[14] 0.01fF
C8252 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# DOUT[6] 0.00fF
C8253 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# DOUT[7] 0.01fF
C8254 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# DOUT[20] 0.00fF
C8255 sky130_fd_sc_hd__dfrtn_1_22/a_651_413# RESET_COUNTERn 0.00fF
C8256 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.00fF
C8257 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_805_47# 0.00fF
C8258 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C8259 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# 0.00fF
C8260 sky130_fd_sc_hd__dfrtn_1_39/a_639_47# VDD 0.01fF
C8261 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_32/a_761_289# 0.01fF
C8262 sky130_fd_sc_hd__inv_1_8/Y sky130_fd_sc_hd__inv_1_8/A 0.08fF
C8263 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# sky130_fd_sc_hd__inv_1_50/Y 0.01fF
C8264 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8265 sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C8266 sky130_fd_sc_hd__inv_1_48/Y DOUT[21] 0.09fF
C8267 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# sky130_fd_sc_hd__dfrtn_1_10/a_543_47# -0.00fF
C8268 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# -0.00fF
C8269 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_3/a_543_47# 0.00fF
C8270 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# 0.00fF
C8271 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__dfrtn_1_3/a_448_47# 0.00fF
C8272 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__dfrtn_1_3/a_805_47# 0.00fF
C8273 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# outb 0.00fF
C8274 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8275 sky130_fd_sc_hd__dfrtn_1_18/a_639_47# VDD 0.00fF
C8276 DOUT[22] DOUT[5] 2.68fF
C8277 sky130_fd_sc_hd__inv_1_38/A sky130_fd_sc_hd__inv_1_38/Y 0.01fF
C8278 sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C8279 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__inv_1_35/Y 0.12fF
C8280 sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# DOUT[2] 0.00fF
C8281 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_448_47# 0.00fF
C8282 sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# sky130_fd_sc_hd__dfrtn_1_19/a_761_289# 0.01fF
C8283 sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C8284 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C8285 sky130_fd_sc_hd__dfrtn_1_16/a_1108_47# RESET_COUNTERn 0.00fF
C8286 sky130_fd_sc_hd__or2_2_0/a_39_297# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C8287 sky130_fd_sc_hd__dfrtn_1_8/a_193_47# RESET_COUNTERn 0.02fF
C8288 sky130_fd_sc_hd__dfrtn_1_8/a_448_47# DOUT[21] 0.00fF
C8289 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# DOUT[14] 0.00fF
C8290 sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8291 VDD sky130_fd_sc_hd__dfrtn_1_9/a_448_47# 0.01fF
C8292 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_20/a_448_47# -0.00fF
C8293 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# -0.00fF
C8294 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C8295 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_805_47# 0.00fF
C8296 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_4/a_1270_413# 0.00fF
C8297 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C8298 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# 0.00fF
C8299 sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C8300 sky130_fd_sc_hd__o2111a_2_0/X sky130_fd_sc_hd__or3_1_0/C 0.00fF
C8301 sky130_fd_sc_hd__o311a_1_0/A3 sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C8302 sky130_fd_sc_hd__o211a_1_1/a_215_47# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C8303 sky130_fd_sc_hd__dfrtn_1_41/a_805_47# sky130_fd_sc_hd__dfrtn_1_38/a_543_47# 0.00fF
C8304 sky130_fd_sc_hd__dfrtn_1_41/a_1270_413# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C8305 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# sky130_fd_sc_hd__dfrtn_1_38/a_805_47# 0.00fF
C8306 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__dfrtn_1_38/a_1270_413# 0.00fF
C8307 sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# sky130_fd_sc_hd__dfrtn_1_38/a_761_289# 0.00fF
C8308 sky130_fd_sc_hd__dfrtn_1_32/a_27_47# sky130_fd_sc_hd__inv_1_36/Y 0.07fF
C8309 sky130_fd_sc_hd__nor3_1_14/a_109_297# DOUT[14] 0.00fF
C8310 sky130_fd_sc_hd__dfrtn_1_19/a_1108_47# VDD 0.07fF
C8311 sky130_fd_sc_hd__dfrtp_1_3/a_1270_413# DOUT[23] 0.00fF
C8312 sky130_fd_sc_hd__nor3_1_10/a_109_297# DOUT[3] 0.00fF
C8313 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__conb_1_0/LO 0.01fF
C8314 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__dfrtn_1_1/a_193_47# 0.00fF
C8315 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# sky130_fd_sc_hd__dfrtn_1_1/a_27_47# 0.00fF
C8316 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_1/a_805_47# 0.00fF
C8317 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# 0.00fF
C8318 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__inv_1_31/A 0.01fF
C8319 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C8320 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__mux4_2_0/a_1281_47# 0.00fF
C8321 sky130_fd_sc_hd__nor3_1_17/a_193_297# VDD 0.00fF
C8322 sky130_fd_sc_hd__or2b_1_0/X sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C8323 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# 0.00fF
C8324 sky130_fd_sc_hd__dfrtn_1_21/a_1462_47# VDD 0.00fF
C8325 sky130_fd_sc_hd__nor3_1_10/a_109_297# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C8326 sky130_fd_sc_hd__dfrtn_1_24/a_805_47# SEL_CONV_TIME[1] 0.00fF
C8327 sky130_fd_sc_hd__dfrtn_1_31/a_543_47# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C8328 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_1217_47# -0.00fF
C8329 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_27/a_761_289# 0.00fF
C8330 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__inv_1_8/Y 0.01fF
C8331 sky130_fd_sc_hd__dfrtn_1_33/a_1462_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C8332 DOUT[4] sky130_fd_sc_hd__dfrtn_1_36/a_761_289# 0.00fF
C8333 sky130_fd_sc_hd__nor3_1_2/a_109_297# VDD 0.00fF
C8334 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C8335 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C8336 sky130_fd_sc_hd__dfrtn_1_23/a_1270_413# RESET_COUNTERn 0.00fF
C8337 sky130_fd_sc_hd__dfrtn_1_22/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8338 sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# sky130_fd_sc_hd__dfrtn_1_26/a_543_47# 0.00fF
C8339 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C8340 sky130_fd_sc_hd__dfrtn_1_10/a_1270_413# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C8341 sky130_fd_sc_hd__dfrtn_1_7/a_651_413# DOUT[6] 0.00fF
C8342 sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# DOUT[20] 0.00fF
C8343 sky130_fd_sc_hd__dfrtn_1_7/a_448_47# DOUT[7] 0.01fF
C8344 sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# RESET_COUNTERn 0.00fF
C8345 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_29/a_543_47# 0.00fF
C8346 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C8347 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.00fF
C8348 sky130_fd_sc_hd__inv_1_0/A DOUT[17] 0.01fF
C8349 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C8350 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_0/a_651_413# -0.00fF
C8351 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# sky130_fd_sc_hd__dfrtn_1_0/a_448_47# -0.00fF
C8352 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# RESET_COUNTERn 0.00fF
C8353 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# DOUT[7] 0.00fF
C8354 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# CLK_REF 0.02fF
C8355 DOUT[7] DOUT[8] 0.04fF
C8356 DOUT[6] RESET_COUNTERn 0.06fF
C8357 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__inv_1_14/A 0.03fF
C8358 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# DOUT[17] 0.00fF
C8359 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# SEL_CONV_TIME[2] 0.00fF
C8360 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_750_97# -0.02fF
C8361 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C8362 sky130_fd_sc_hd__dfrtn_1_26/a_761_289# sky130_fd_sc_hd__dfrtn_1_27/a_448_47# 0.00fF
C8363 sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# sky130_fd_sc_hd__dfrtn_1_27/a_543_47# 0.00fF
C8364 sky130_fd_sc_hd__dfrtn_1_26/a_651_413# sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.00fF
C8365 sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C8366 sky130_fd_sc_hd__nor3_1_9/a_109_297# DOUT[3] 0.00fF
C8367 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__o311a_1_0/a_266_47# 0.00fF
C8368 sky130_fd_sc_hd__dfrtn_1_24/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8369 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# VDD 0.00fF
C8370 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C8371 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__inv_1_33/A 0.01fF
C8372 CLK_REF sky130_fd_sc_hd__dfrtn_1_21/a_27_47# 0.01fF
C8373 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# 0.00fF
C8374 sky130_fd_sc_hd__dfrtn_1_16/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8375 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8376 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# VDD 0.07fF
C8377 sky130_fd_sc_hd__dfrtn_1_11/a_1462_47# outb 0.00fF
C8378 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__dfrtn_1_3/a_651_413# 0.00fF
C8379 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__inv_1_53/A 0.01fF
C8380 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C8381 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C8382 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_31/a_1283_21# 0.00fF
C8383 sky130_fd_sc_hd__nor3_2_0/A sky130_fd_sc_hd__inv_1_1/A 0.00fF
C8384 sky130_fd_sc_hd__inv_1_6/A DOUT[3] 0.02fF
C8385 sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# DOUT[14] 0.00fF
C8386 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_12/a_27_47# 0.02fF
C8387 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__or2_2_0/A 0.26fF
C8388 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__mux4_2_0/a_872_316# 0.00fF
C8389 sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# sky130_fd_sc_hd__dfrtn_1_19/a_448_47# 0.00fF
C8390 sky130_fd_sc_hd__inv_1_1/A DOUT[17] 0.03fF
C8391 sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C8392 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.01fF
C8393 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C8394 sky130_fd_sc_hd__dfrtn_1_8/a_1462_47# RESET_COUNTERn 0.00fF
C8395 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_14/a_27_47# 0.00fF
C8396 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_14/a_193_47# 0.00fF
C8397 sky130_fd_sc_hd__dfrtp_1_0/a_1270_413# sky130_fd_sc_hd__o211a_1_0/X 0.00fF
C8398 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_6/A 0.76fF
C8399 sky130_fd_sc_hd__dfrtn_1_30/a_639_47# SEL_CONV_TIME[1] 0.00fF
C8400 sky130_fd_sc_hd__dfrtn_1_20/a_805_47# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C8401 sky130_fd_sc_hd__o211a_1_0/X out 0.00fF
C8402 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_13/A 0.01fF
C8403 sky130_fd_sc_hd__dfrtn_1_23/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8404 sky130_fd_sc_hd__or3b_2_0/a_388_297# sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# 0.00fF
C8405 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# VDD 0.11fF
C8406 sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C8407 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_18/a_761_289# 0.00fF
C8408 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__o221ai_1_0/a_295_297# 0.00fF
C8409 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8410 sky130_fd_sc_hd__nand3b_1_1/a_232_47# SEL_CONV_TIME[0] 0.00fF
C8411 sky130_fd_sc_hd__or3_1_0/a_111_297# SEL_CONV_TIME[0] 0.00fF
C8412 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C8413 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__nor3_1_3/a_193_297# 0.00fF
C8414 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8415 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# VDD 0.08fF
C8416 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_44/A 0.01fF
C8417 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C8418 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C8419 sky130_fd_sc_hd__dfrtn_1_38/a_761_289# SEL_CONV_TIME[1] 0.00fF
C8420 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# RESET_COUNTERn 0.06fF
C8421 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8422 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__dfrtn_1_30/a_193_47# 0.00fF
C8423 sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C8424 sky130_fd_sc_hd__nor3_2_3/B DOUT[21] 0.46fF
C8425 sky130_fd_sc_hd__nor3_1_10/a_109_297# DOUT[20] 0.00fF
C8426 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C8427 sky130_fd_sc_hd__dfrtn_1_33/a_543_47# VDD 0.05fF
C8428 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__inv_1_27/Y 0.00fF
C8429 sky130_fd_sc_hd__dfrtn_1_30/a_1270_413# VDD 0.00fF
C8430 sky130_fd_sc_hd__dfrtn_1_31/a_761_289# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C8431 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# DOUT[3] 0.00fF
C8432 sky130_fd_sc_hd__mux4_2_0/a_600_345# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C8433 sky130_fd_sc_hd__nand2_1_2/Y SEL_CONV_TIME[0] 0.15fF
C8434 sky130_fd_sc_hd__dfrtn_1_4/a_805_47# DOUT[3] 0.00fF
C8435 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C8436 sky130_fd_sc_hd__inv_1_29/A RESET_COUNTERn 0.70fF
C8437 sky130_fd_sc_hd__dfrtn_1_20/a_543_47# sky130_fd_sc_hd__inv_1_35/A 0.01fF
C8438 sky130_fd_sc_hd__dfrtn_1_16/a_1270_413# DOUT[23] 0.00fF
C8439 sky130_fd_sc_hd__or3b_2_0/B RESET_COUNTERn 0.25fF
C8440 DOUT[4] sky130_fd_sc_hd__dfrtn_1_31/a_1283_21# 0.00fF
C8441 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__inv_1_41/Y 0.01fF
C8442 sky130_fd_sc_hd__dfrtn_1_30/a_651_413# sky130_fd_sc_hd__dfrtn_1_31/a_27_47# 0.00fF
C8443 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__dfrtn_1_31/a_448_47# 0.00fF
C8444 sky130_fd_sc_hd__dfrtn_1_30/a_448_47# sky130_fd_sc_hd__dfrtn_1_31/a_193_47# 0.00fF
C8445 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_651_413# 0.00fF
C8446 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C8447 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# DOUT[14] 0.00fF
C8448 sky130_fd_sc_hd__dfrtn_1_14/a_639_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C8449 sky130_fd_sc_hd__dfrtn_1_35/a_193_47# sky130_fd_sc_hd__dfrtn_1_35/a_639_47# -0.00fF
C8450 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C8451 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# SEL_CONV_TIME[1] 0.00fF
C8452 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# 0.00fF
C8453 sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# DOUT[17] 0.00fF
C8454 sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# SEL_CONV_TIME[1] 0.00fF
C8455 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__dfrtn_1_17/a_448_47# 0.00fF
C8456 sky130_fd_sc_hd__o211a_1_1/a_510_47# sky130_fd_sc_hd__dfrtn_1_17/a_543_47# 0.00fF
C8457 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C8458 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_543_47# 0.00fF
C8459 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C8460 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_29/a_761_289# 0.00fF
C8461 sky130_fd_sc_hd__dfrtn_1_25/a_651_413# SEL_CONV_TIME[0] 0.00fF
C8462 sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__o211a_1_0/a_510_47# 0.00fF
C8463 sky130_fd_sc_hd__nor3_1_7/a_193_297# DOUT[19] 0.00fF
C8464 sky130_fd_sc_hd__nand3b_1_1/a_53_93# DOUT[21] 0.01fF
C8465 sky130_fd_sc_hd__o311a_1_0/A3 sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C8466 sky130_fd_sc_hd__or3_1_0/a_29_53# DOUT[21] 0.00fF
C8467 sky130_fd_sc_hd__dfrtn_1_38/a_193_47# VDD 0.14fF
C8468 sky130_fd_sc_hd__dfrtn_1_36/a_805_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C8469 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__dfrtn_1_11/a_193_47# 0.00fF
C8470 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# 0.00fF
C8471 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# 0.00fF
C8472 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# sky130_fd_sc_hd__dfrtn_1_11/a_27_47# 0.00fF
C8473 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_11/a_448_47# 0.00fF
C8474 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_651_413# 0.00fF
C8475 sky130_fd_sc_hd__o211a_1_1/a_510_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8476 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C8477 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C8478 sky130_fd_sc_hd__inv_1_36/A sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C8479 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_12/a_1217_47# 0.00fF
C8480 DOUT[4] sky130_fd_sc_hd__dfrtn_1_32/a_639_47# 0.00fF
C8481 DOUT[9] sky130_fd_sc_hd__nor3_1_3/a_193_297# -0.00fF
C8482 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/a_543_47# -0.00fF
C8483 sky130_fd_sc_hd__dfrtn_1_7/a_543_47# sky130_fd_sc_hd__inv_1_6/A 0.01fF
C8484 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# 0.00fF
C8485 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__dfrtn_1_40/a_651_413# 0.00fF
C8486 sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C8487 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_17/a_1270_413# 0.00fF
C8488 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__dfrtn_1_17/a_639_47# 0.00fF
C8489 sky130_fd_sc_hd__dfrtp_1_2/a_639_47# sky130_fd_sc_hd__dfrtn_1_17/a_543_47# 0.00fF
C8490 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_17/a_805_47# 0.00fF
C8491 sky130_fd_sc_hd__dfrtp_1_2/a_448_47# sky130_fd_sc_hd__dfrtn_1_17/a_448_47# 0.00fF
C8492 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# 0.00fF
C8493 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# 0.00fF
C8494 sky130_fd_sc_hd__dfrtn_1_12/a_651_413# sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# 0.00fF
C8495 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C8496 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__dfrtn_1_37/a_761_289# -0.00fF
C8497 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_37/a_543_47# -0.00fF
C8498 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_14/a_448_47# 0.00fF
C8499 sky130_fd_sc_hd__dfrtn_1_28/a_1283_21# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C8500 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8501 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__dfrtn_1_42/a_639_47# 0.00fF
C8502 sky130_fd_sc_hd__dfrtn_1_26/a_543_47# VDD 0.04fF
C8503 sky130_fd_sc_hd__o211a_1_0/a_510_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C8504 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C8505 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# DOUT[14] 0.00fF
C8506 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C8507 sky130_fd_sc_hd__nor3_1_3/a_109_297# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C8508 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C8509 sky130_fd_sc_hd__nor3_2_0/a_281_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8510 sky130_fd_sc_hd__inv_1_6/A DOUT[20] 0.08fF
C8511 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_41/Y 0.19fF
C8512 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8513 sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# VDD 0.10fF
C8514 DOUT[4] sky130_fd_sc_hd__or2b_1_0/a_27_53# 0.00fF
C8515 sky130_fd_sc_hd__dfrtp_1_2/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8516 DOUT[4] sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C8517 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_7/a_193_47# 0.00fF
C8518 sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# VDD 0.00fF
C8519 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# 0.00fF
C8520 sky130_fd_sc_hd__or2b_1_0/a_301_297# sky130_fd_sc_hd__dfrtn_1_30/a_761_289# 0.00fF
C8521 sky130_fd_sc_hd__dfrtn_1_23/a_543_47# sky130_fd_sc_hd__inv_1_40/Y 0.02fF
C8522 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_193_47# -0.29fF
C8523 sky130_fd_sc_hd__dfrtn_1_28/a_1283_21# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C8524 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C8525 DOUT[23] RESET_COUNTERn 0.03fF
C8526 sky130_fd_sc_hd__dfrtn_1_16/a_651_413# sky130_fd_sc_hd__inv_1_26/A 0.00fF
C8527 sky130_fd_sc_hd__o2111a_2_0/a_674_297# SEL_CONV_TIME[1] 0.00fF
C8528 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# RESET_COUNTERn 0.01fF
C8529 sky130_fd_sc_hd__dfrtn_1_25/a_448_47# DOUT[21] 0.00fF
C8530 sky130_fd_sc_hd__dfrtn_1_42/a_1462_47# sky130_fd_sc_hd__dfrtn_1_23/a_193_47# 0.00fF
C8531 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_6/a_651_413# 0.00fF
C8532 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C8533 sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# RESET_COUNTERn 0.00fF
C8534 sky130_fd_sc_hd__nor3_1_4/a_109_297# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C8535 sky130_fd_sc_hd__dfrtn_1_32/a_448_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C8536 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__inv_1_13/Y 0.01fF
C8537 sky130_fd_sc_hd__dfrtn_1_33/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8538 sky130_fd_sc_hd__nor3_1_19/a_109_297# SEL_CONV_TIME[1] 0.00fF
C8539 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# DOUT[15] 0.00fF
C8540 sky130_fd_sc_hd__dfrtn_1_3/a_805_47# RESET_COUNTERn 0.00fF
C8541 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__inv_1_49/A 0.01fF
C8542 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__inv_1_43/A 0.01fF
C8543 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__dfrtn_1_9/a_448_47# 0.00fF
C8544 sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# HEADER_0/a_508_138# 0.00fF
C8545 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8546 sky130_fd_sc_hd__nand2_1_1/Y DOUT[21] 0.00fF
C8547 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# VDD 0.01fF
C8548 sky130_fd_sc_hd__dfrtn_1_42/a_761_289# RESET_COUNTERn 0.02fF
C8549 sky130_fd_sc_hd__mux4_2_0/a_288_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C8550 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# SEL_CONV_TIME[3] 0.00fF
C8551 sky130_fd_sc_hd__dfrtn_1_34/a_448_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C8552 sky130_fd_sc_hd__dfrtn_1_21/a_448_47# sky130_fd_sc_hd__inv_1_35/A 0.00fF
C8553 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C8554 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_10/a_761_289# 0.00fF
C8555 sky130_fd_sc_hd__dfrtn_1_0/a_448_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C8556 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C8557 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_543_47# 0.00fF
C8558 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C8559 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C8560 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# HEADER_0/a_508_138# 0.00fF
C8561 sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C8562 HEADER_0/a_508_138# DOUT[6] 0.00fF
C8563 sky130_fd_sc_hd__dfrtn_1_0/a_639_47# DOUT[17] 0.00fF
C8564 sky130_fd_sc_hd__o2111a_2_0/a_80_21# VDD 0.09fF
C8565 DOUT[13] sky130_fd_sc_hd__dfrtn_1_36/a_1270_413# 0.00fF
C8566 sky130_fd_sc_hd__dfrtn_1_24/a_651_413# sky130_fd_sc_hd__dfrtn_1_29/a_651_413# 0.00fF
C8567 sky130_fd_sc_hd__dfrtn_1_17/a_448_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C8568 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# DOUT[6] 0.00fF
C8569 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# DOUT[20] 0.00fF
C8570 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# RESET_COUNTERn 0.02fF
C8571 sky130_fd_sc_hd__dfrtn_1_4/a_448_47# RESET_COUNTERn 0.01fF
C8572 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# SEL_CONV_TIME[0] 0.00fF
C8573 sky130_fd_sc_hd__dfrtn_1_38/a_1462_47# VDD 0.00fF
C8574 sky130_fd_sc_hd__dfrtn_1_33/a_805_47# sky130_fd_sc_hd__inv_1_45/A 0.00fF
C8575 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_49/A 0.04fF
C8576 sky130_fd_sc_hd__dfrtp_1_1/D sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C8577 DOUT[15] sky130_fd_sc_hd__inv_1_40/Y 0.01fF
C8578 DOUT[13] VDD 2.51fF
C8579 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__dfrtn_1_34/a_27_47# 0.00fF
C8580 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__dfrtn_1_11/a_1462_47# 0.00fF
C8581 sky130_fd_sc_hd__dfrtn_1_42/a_805_47# DOUT[15] 0.00fF
C8582 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# sky130_fd_sc_hd__inv_1_49/A 0.25fF
C8583 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__o311a_1_0/A3 0.02fF
C8584 DOUT[1] sky130_fd_sc_hd__inv_1_37/A 0.02fF
C8585 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.01fF
C8586 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# SEL_CONV_TIME[2] 0.02fF
C8587 VDD sky130_fd_sc_hd__inv_1_8/A 0.56fF
C8588 CLK_REF sky130_fd_sc_hd__or2_2_0/A 0.13fF
C8589 sky130_fd_sc_hd__dfrtn_1_14/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8590 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# VDD 0.08fF
C8591 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# 0.00fF
C8592 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# 0.00fF
C8593 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C8594 sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8595 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# DOUT[3] 0.00fF
C8596 sky130_fd_sc_hd__dfrtp_1_0/a_1283_21# RESET_COUNTERn 0.03fF
C8597 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C8598 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__dfrtn_1_41/a_651_413# -0.00fF
C8599 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C8600 sky130_fd_sc_hd__o2111a_2_0/a_386_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C8601 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_38/a_1270_413# 0.00fF
C8602 sky130_fd_sc_hd__dfrtn_1_3/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8603 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_8/a_639_47# 0.00fF
C8604 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# sky130_fd_sc_hd__inv_1_2/Y 0.01fF
C8605 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C8606 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__nor3_1_5/a_193_297# 0.00fF
C8607 sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# RESET_COUNTERn 0.01fF
C8608 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C8609 sky130_fd_sc_hd__dfrtn_1_22/a_543_47# sky130_fd_sc_hd__inv_1_39/Y 0.01fF
C8610 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_13/A 0.63fF
C8611 sky130_fd_sc_hd__dfrtn_1_25/a_1462_47# RESET_COUNTERn 0.00fF
C8612 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.03fF
C8613 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C8614 sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C8615 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C8616 sky130_fd_sc_hd__inv_1_31/A RESET_COUNTERn 0.57fF
C8617 sky130_fd_sc_hd__dfrtp_1_3/a_448_47# sky130_fd_sc_hd__o211a_1_1/a_510_47# 0.00fF
C8618 sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# RESET_COUNTERn 0.01fF
C8619 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8620 sky130_fd_sc_hd__dfrtp_1_0/a_1462_47# DOUT[15] 0.00fF
C8621 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_26/a_805_47# 0.00fF
C8622 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C8623 sky130_fd_sc_hd__nor3_1_10/a_193_297# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C8624 sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C8625 en DOUT[8] 0.03fF
C8626 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# SEL_CONV_TIME[3] 0.00fF
C8627 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_1270_413# 0.00fF
C8628 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C8629 sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# SEL_CONV_TIME[3] 0.00fF
C8630 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__nor3_2_0/a_27_297# 0.01fF
C8631 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# DOUT[3] 0.00fF
C8632 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# VDD 0.16fF
C8633 sky130_fd_sc_hd__mux4_2_0/a_872_316# sky130_fd_sc_hd__o311a_1_0/a_266_47# 0.00fF
C8634 sky130_fd_sc_hd__dfrtn_1_9/a_761_289# RESET_COUNTERn 0.02fF
C8635 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtp_1_3/a_805_47# 0.00fF
C8636 sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# sky130_fd_sc_hd__dfrtp_1_3/a_543_47# 0.00fF
C8637 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# sky130_fd_sc_hd__dfrtp_1_3/a_651_413# 0.00fF
C8638 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__mux4_2_0/a_872_316# -0.00fF
C8639 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C8640 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# 0.00fF
C8641 sky130_fd_sc_hd__inv_1_45/Y sky130_fd_sc_hd__inv_1_43/A 0.01fF
C8642 sky130_fd_sc_hd__dfrtn_1_19/a_193_47# RESET_COUNTERn 0.00fF
C8643 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C8644 CLK_REF sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# 0.00fF
C8645 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__inv_1_2/A 0.01fF
C8646 sky130_fd_sc_hd__mux4_2_0/a_288_47# sky130_fd_sc_hd__inv_1_32/A 0.01fF
C8647 sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# SEL_CONV_TIME[0] 0.00fF
C8648 sky130_fd_sc_hd__o221ai_1_0/a_109_47# RESET_COUNTERn 0.00fF
C8649 sky130_fd_sc_hd__or3_1_0/a_183_297# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C8650 sky130_fd_sc_hd__inv_1_0/Y DOUT[18] 0.01fF
C8651 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__o2111a_2_0/a_458_47# 0.00fF
C8652 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_3/A 0.00fF
C8653 sky130_fd_sc_hd__dfrtp_1_0/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8654 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C8655 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C8656 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__inv_1_8/A 0.32fF
C8657 sky130_fd_sc_hd__inv_1_18/Y VIN 0.34fF
C8658 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C8659 sky130_fd_sc_hd__inv_1_33/A RESET_COUNTERn 0.15fF
C8660 sky130_fd_sc_hd__nor3_2_1/a_281_297# sky130_fd_sc_hd__conb_1_0/LO 0.00fF
C8661 sky130_fd_sc_hd__dfrtn_1_31/a_1462_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C8662 sky130_fd_sc_hd__dfrtn_1_35/a_1283_21# DOUT[16] 0.00fF
C8663 sky130_fd_sc_hd__dfrtn_1_35/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.00fF
C8664 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# 0.00fF
C8665 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# -0.00fF
C8666 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# -0.00fF
C8667 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# sky130_fd_sc_hd__dfrtn_1_25/a_543_47# -0.00fF
C8668 DOUT[13] sky130_fd_sc_hd__dfrtn_1_31/a_805_47# 0.00fF
C8669 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# 0.00fF
C8670 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_1270_413# 0.00fF
C8671 sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# SEL_CONV_TIME[2] 0.00fF
C8672 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_29/a_805_47# 0.00fF
C8673 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C8674 sky130_fd_sc_hd__dfrtn_1_28/a_1270_413# VDD 0.00fF
C8675 sky130_fd_sc_hd__dfrtn_1_29/a_639_47# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C8676 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C8677 sky130_fd_sc_hd__dfrtn_1_4/a_448_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C8678 sky130_fd_sc_hd__dfrtn_1_25/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8679 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__nor3_2_0/A 0.01fF
C8680 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_37/a_543_47# 0.02fF
C8681 sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# sky130_fd_sc_hd__inv_1_12/A 0.02fF
C8682 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# VDD 0.08fF
C8683 sky130_fd_sc_hd__dfrtn_1_16/a_1108_47# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C8684 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__inv_1_14/A 0.01fF
C8685 VDD sky130_fd_sc_hd__inv_1_27/Y 0.15fF
C8686 sky130_fd_sc_hd__mux4_1_0/a_1478_413# SEL_CONV_TIME[1] 0.00fF
C8687 DOUT[9] sky130_fd_sc_hd__nor3_2_3/B 1.08fF
C8688 sky130_fd_sc_hd__nor3_1_10/a_193_297# DOUT[9] 0.00fF
C8689 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C8690 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.01fF
C8691 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C8692 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_14/a_27_47# 0.02fF
C8693 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__nor3_2_3/C 0.37fF
C8694 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__inv_1_6/A 0.01fF
C8695 sky130_fd_sc_hd__dfrtn_1_39/a_761_289# sky130_fd_sc_hd__inv_1_32/Y 0.00fF
C8696 sky130_fd_sc_hd__dfrtn_1_20/a_448_47# VDD 0.01fF
C8697 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C8698 sky130_fd_sc_hd__dfrtn_1_24/a_805_47# DOUT[21] 0.00fF
C8699 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# RESET_COUNTERn 0.00fF
C8700 sky130_fd_sc_hd__dfrtn_1_42/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8701 sky130_fd_sc_hd__dfrtn_1_25/a_1270_413# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C8702 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# RESET_COUNTERn 0.05fF
C8703 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C8704 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C8705 sky130_fd_sc_hd__nor3_1_10/a_109_297# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C8706 DOUT[1] sky130_fd_sc_hd__dfrtn_1_36/a_448_47# 0.00fF
C8707 DOUT[4] sky130_fd_sc_hd__dfrtn_1_8/a_1108_47# 0.00fF
C8708 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.01fF
C8709 sky130_fd_sc_hd__dfrtn_1_20/a_639_47# sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# 0.00fF
C8710 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_4/a_543_47# 0.00fF
C8711 sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__inv_1_23/A 0.00fF
C8712 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8713 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_26/a_651_413# 0.00fF
C8714 sky130_fd_sc_hd__or3_1_0/C sky130_fd_sc_hd__inv_1_43/A 0.02fF
C8715 sky130_fd_sc_hd__dfrtn_1_16/a_543_47# DOUT[2] 0.01fF
C8716 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# sky130_fd_sc_hd__dfrtn_1_42/a_651_413# -0.00fF
C8717 sky130_fd_sc_hd__dfrtn_1_42/a_193_47# sky130_fd_sc_hd__dfrtn_1_42/a_448_47# -0.00fF
C8718 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_27_47# 0.00fF
C8719 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_193_47# 0.00fF
C8720 sky130_fd_sc_hd__o221ai_1_0/a_295_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8721 HEADER_2/a_508_138# DOUT[11] 0.02fF
C8722 DOUT[9] sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C8723 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# DOUT[11] 0.00fF
C8724 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__mux4_1_0/X 0.01fF
C8725 sky130_fd_sc_hd__dfrtn_1_30/a_805_47# SEL_CONV_TIME[0] 0.00fF
C8726 sky130_fd_sc_hd__nor3_1_4/a_193_297# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C8727 sky130_fd_sc_hd__dfrtp_1_1/D DOUT[0] 0.00fF
C8728 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8729 sky130_fd_sc_hd__inv_1_31/A SEL_CONV_TIME[3] 0.02fF
C8730 sky130_fd_sc_hd__mux4_1_0/a_1290_413# VDD 0.09fF
C8731 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C8732 sky130_fd_sc_hd__dfrtn_1_10/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8733 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C8734 sky130_fd_sc_hd__dfrtn_1_10/a_1217_47# VDD 0.00fF
C8735 sky130_fd_sc_hd__o211a_1_0/a_79_21# VDD 0.08fF
C8736 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# VIN 0.09fF
C8737 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# 0.00fF
C8738 sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C8739 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# sky130_fd_sc_hd__dfrtn_1_15/a_543_47# 0.00fF
C8740 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# DOUT[23] 0.00fF
C8741 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_20/a_761_289# 0.00fF
C8742 sky130_fd_sc_hd__dfrtn_1_24/a_805_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C8743 DOUT[23] DOUT[10] 0.03fF
C8744 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C8745 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# -0.00fF
C8746 sky130_fd_sc_hd__dfrtn_1_27/a_761_289# sky130_fd_sc_hd__dfrtn_1_27/a_543_47# -0.00fF
C8747 sky130_fd_sc_hd__nor3_1_9/a_193_297# DOUT[9] 0.00fF
C8748 sky130_fd_sc_hd__dfrtn_1_19/a_1462_47# RESET_COUNTERn 0.00fF
C8749 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C8750 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# 0.00fF
C8751 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C8752 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C8753 sky130_fd_sc_hd__mux4_2_0/a_1060_369# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C8754 sky130_fd_sc_hd__dfrtn_1_38/a_543_47# SEL_CONV_TIME[0] 0.00fF
C8755 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_639_47# -0.00fF
C8756 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# DOUT[20] 0.00fF
C8757 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# RESET_COUNTERn 0.04fF
C8758 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__inv_1_8/A 0.00fF
C8759 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_4/a_805_47# 0.00fF
C8760 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_4/a_1270_413# 0.00fF
C8761 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C8762 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C8763 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_4/a_651_413# 0.00fF
C8764 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_761_289# -0.00fF
C8765 sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C8766 sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# SEL_CONV_TIME[2] 0.01fF
C8767 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C8768 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C8769 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__o311a_1_0/a_368_297# 0.00fF
C8770 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.00fF
C8771 sky130_fd_sc_hd__inv_1_31/A SEL_CONV_TIME[2] 0.03fF
C8772 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__o311a_1_0/a_266_297# 0.00fF
C8773 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# 0.00fF
C8774 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__inv_1_45/A 0.06fF
C8775 sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# SEL_CONV_TIME[2] 0.00fF
C8776 sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# DOUT[21] 0.00fF
C8777 DOUT[1] sky130_fd_sc_hd__dfrtn_1_32/a_761_289# 0.00fF
C8778 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C8779 sky130_fd_sc_hd__dfrtn_1_27/a_639_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C8780 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.00fF
C8781 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__mux4_2_0/a_372_413# 0.00fF
C8782 sky130_fd_sc_hd__dfrtn_1_12/a_1217_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C8783 sky130_fd_sc_hd__dfrtn_1_0/a_1462_47# VDD 0.00fF
C8784 sky130_fd_sc_hd__dfrtn_1_35/a_1270_413# VDD 0.00fF
C8785 sky130_fd_sc_hd__o311a_1_0/a_266_47# SEL_CONV_TIME[1] 0.00fF
C8786 sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# RESET_COUNTERn 0.01fF
C8787 sky130_fd_sc_hd__dfrtn_1_12/a_1270_413# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C8788 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.00fF
C8789 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C8790 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_6/Y 0.27fF
C8791 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_6/A 0.01fF
C8792 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C8793 sky130_fd_sc_hd__dfrtn_1_18/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_761_289# -0.00fF
C8794 sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# SEL_CONV_TIME[0] 0.01fF
C8795 sky130_fd_sc_hd__dfrtn_1_3/a_1462_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C8796 sky130_fd_sc_hd__mux4_2_0/a_788_316# SEL_CONV_TIME[1] 0.05fF
C8797 sky130_fd_sc_hd__inv_1_33/A SEL_CONV_TIME[3] 0.06fF
C8798 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# DOUT[19] 0.01fF
C8799 sky130_fd_sc_hd__dfrtn_1_27/a_651_413# sky130_fd_sc_hd__or3_1_0/C 0.01fF
C8800 sky130_fd_sc_hd__dfrtn_1_34/a_448_47# SEL_CONV_TIME[0] 0.00fF
C8801 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C8802 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# VDD 0.07fF
C8803 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# 0.00fF
C8804 sky130_fd_sc_hd__dfrtn_1_23/a_639_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C8805 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_30/a_448_47# 0.00fF
C8806 sky130_fd_sc_hd__inv_1_0/Y DOUT[22] 0.00fF
C8807 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C8808 sky130_fd_sc_hd__dfrtn_1_30/a_761_289# DONE 0.00fF
C8809 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_639_47# -0.00fF
C8810 sky130_fd_sc_hd__dfrtp_1_0/a_1283_21# SLC_0/a_264_22# 0.00fF
C8811 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# sky130_fd_sc_hd__inv_1_25/A 0.00fF
C8812 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# RESET_COUNTERn 0.00fF
C8813 sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C8814 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# sky130_fd_sc_hd__inv_1_26/A 0.00fF
C8815 sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8816 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__nand3b_1_0/a_232_47# 0.00fF
C8817 sky130_fd_sc_hd__dfrtn_1_41/a_1270_413# SEL_CONV_TIME[1] 0.00fF
C8818 sky130_fd_sc_hd__or2_2_0/X RESET_COUNTERn 0.03fF
C8819 CLK_REF sky130_fd_sc_hd__dfrtp_1_3/a_1270_413# 0.00fF
C8820 DOUT[1] DOUT[14] 0.00fF
C8821 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# 0.00fF
C8822 sky130_fd_sc_hd__dfrtn_1_8/a_1108_47# outb 0.00fF
C8823 sky130_fd_sc_hd__o211a_1_1/a_297_297# RESET_COUNTERn 0.00fF
C8824 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8825 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_12/a_1217_47# -0.00fF
C8826 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_10/a_27_47# 0.26fF
C8827 sky130_fd_sc_hd__dfrtn_1_10/a_1270_413# sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# 0.00fF
C8828 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# 0.00fF
C8829 DOUT[9] sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# 0.00fF
C8830 sky130_fd_sc_hd__dfrtn_1_7/a_448_47# VIN 0.01fF
C8831 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_6/Y 0.20fF
C8832 sky130_fd_sc_hd__o311a_1_0/a_81_21# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C8833 sky130_fd_sc_hd__o311a_1_0/a_368_297# VDD 0.00fF
C8834 sky130_fd_sc_hd__inv_1_33/A SEL_CONV_TIME[2] 0.29fF
C8835 sky130_fd_sc_hd__dfrtn_1_21/a_1270_413# sky130_fd_sc_hd__inv_1_35/Y 0.00fF
C8836 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# 0.00fF
C8837 DOUT[9] sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# 0.00fF
C8838 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# DOUT[11] 0.00fF
C8839 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__inv_1_5/Y -0.02fF
C8840 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# SEL_CONV_TIME[3] 0.00fF
C8841 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C8842 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# DOUT[5] 0.00fF
C8843 sky130_fd_sc_hd__o2111a_2_0/X RESET_COUNTERn 0.00fF
C8844 sky130_fd_sc_hd__mux4_2_0/a_372_413# VDD 0.01fF
C8845 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# out 0.01fF
C8846 sky130_fd_sc_hd__or2_2_0/a_121_297# VDD 0.00fF
C8847 sky130_fd_sc_hd__inv_1_4/Y DOUT[6] 0.08fF
C8848 sky130_fd_sc_hd__dfrtn_1_27/a_193_47# SEL_CONV_TIME[1] 0.00fF
C8849 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# VIN 0.00fF
C8850 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__inv_1_53/A 0.01fF
C8851 VIN DOUT[8] 2.70fF
C8852 sky130_fd_sc_hd__mux4_2_0/X RESET_COUNTERn 0.00fF
C8853 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__nor3_2_1/a_281_297# 0.00fF
C8854 VDD sky130_fd_sc_hd__nor3_1_4/A 0.58fF
C8855 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__inv_1_43/Y 0.01fF
C8856 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C8857 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__nand3b_1_1/Y -0.00fF
C8858 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__nand2_1_1/a_113_47# 0.00fF
C8859 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C8860 sky130_fd_sc_hd__o2111a_2_0/a_386_47# SEL_CONV_TIME[0] 0.00fF
C8861 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# RESET_COUNTERn 0.01fF
C8862 sky130_fd_sc_hd__dfrtn_1_35/a_543_47# sky130_fd_sc_hd__inv_1_38/Y 0.01fF
C8863 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C8864 sky130_fd_sc_hd__dfrtn_1_11/a_761_289# VDD 0.05fF
C8865 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# RESET_COUNTERn 0.00fF
C8866 sky130_fd_sc_hd__dfrtn_1_35/a_761_289# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C8867 sky130_fd_sc_hd__inv_1_45/Y sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8868 sky130_fd_sc_hd__nor3_1_20/a_109_297# VDD 0.00fF
C8869 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8870 sky130_fd_sc_hd__dfrtn_1_30/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8871 sky130_fd_sc_hd__dfrtn_1_41/a_651_413# VDD 0.01fF
C8872 sky130_fd_sc_hd__nor3_1_4/a_193_297# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C8873 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C8874 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# RESET_COUNTERn 0.00fF
C8875 sky130_fd_sc_hd__nor3_1_19/a_193_297# SEL_CONV_TIME[0] 0.00fF
C8876 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_34/a_761_289# 0.00fF
C8877 sky130_fd_sc_hd__dfrtn_1_8/a_27_47# sky130_fd_sc_hd__inv_1_8/A 0.02fF
C8878 sky130_fd_sc_hd__nand3b_1_0/a_316_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8879 sky130_fd_sc_hd__dfrtn_1_21/a_193_47# sky130_fd_sc_hd__dfrtn_1_19/a_1108_47# 0.00fF
C8880 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_39/a_1270_413# 0.00fF
C8881 sky130_fd_sc_hd__o311a_1_0/a_585_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C8882 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__mux4_1_0/a_27_413# 0.00fF
C8883 sky130_fd_sc_hd__dfrtn_1_39/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_1462_47# 0.00fF
C8884 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__dfrtn_1_14/a_651_413# 0.00fF
C8885 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_30/a_651_413# 0.00fF
C8886 sky130_fd_sc_hd__dfrtn_1_33/a_805_47# RESET_COUNTERn 0.00fF
C8887 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__mux4_2_0/a_1281_47# 0.00fF
C8888 sky130_fd_sc_hd__mux4_2_0/a_600_345# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C8889 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8890 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_18/a_1270_413# 0.00fF
C8891 VDD sky130_fd_sc_hd__inv_1_15/A 2.05fF
C8892 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C8893 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C8894 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# VDD 0.16fF
C8895 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# 0.00fF
C8896 sky130_fd_sc_hd__dfrtn_1_3/a_639_47# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.00fF
C8897 sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C8898 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.05fF
C8899 sky130_fd_sc_hd__o211a_1_0/a_79_21# sky130_fd_sc_hd__o211a_1_0/X 0.01fF
C8900 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# RESET_COUNTERn 0.03fF
C8901 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/D 0.00fF
C8902 sky130_fd_sc_hd__dfrtn_1_21/a_543_47# RESET_COUNTERn 0.02fF
C8903 sky130_fd_sc_hd__dfrtn_1_37/a_1270_413# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C8904 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C8905 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C8906 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C8907 sky130_fd_sc_hd__nand2_1_1/a_113_47# VDD 0.00fF
C8908 sky130_fd_sc_hd__o2111a_2_0/a_674_297# DOUT[21] 0.00fF
C8909 sky130_fd_sc_hd__nor3_2_2/A DOUT[23] 0.00fF
C8910 sky130_fd_sc_hd__inv_1_25/A DOUT[15] 0.04fF
C8911 sky130_fd_sc_hd__o221ai_1_0/a_493_297# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C8912 sky130_fd_sc_hd__dfrtn_1_16/a_1217_47# sky130_fd_sc_hd__inv_1_25/A 0.00fF
C8913 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C8914 sky130_fd_sc_hd__dfrtn_1_38/a_1270_413# RESET_COUNTERn 0.00fF
C8915 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__inv_1_43/Y 0.03fF
C8916 sky130_fd_sc_hd__dfrtn_1_14/a_805_47# DOUT[18] 0.00fF
C8917 CLK_REF sky130_fd_sc_hd__dfrtn_1_21/a_1270_413# 0.00fF
C8918 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8919 sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C8920 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# VDD 0.04fF
C8921 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C8922 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C8923 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C8924 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_448_47# 0.00fF
C8925 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.00fF
C8926 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_36/Y 0.03fF
C8927 sky130_fd_sc_hd__nor3_1_19/a_109_297# DOUT[21] 0.00fF
C8928 sky130_fd_sc_hd__dfrtp_1_3/a_761_289# sky130_fd_sc_hd__or2_2_0/B 0.02fF
C8929 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8930 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# VDD 0.06fF
C8931 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_30/a_193_47# 0.00fF
C8932 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_10/a_1217_47# 0.00fF
C8933 sky130_fd_sc_hd__dfrtn_1_39/a_1270_413# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C8934 sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C8935 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__or3_1_0/C 0.01fF
C8936 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__inv_1_49/A 0.01fF
C8937 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8938 sky130_fd_sc_hd__mux4_2_0/a_1281_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8939 sky130_fd_sc_hd__dfrtn_1_33/a_761_289# DOUT[23] 0.00fF
C8940 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# DOUT[5] 0.00fF
C8941 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_448_47# -0.00fF
C8942 sky130_fd_sc_hd__dfrtn_1_9/a_448_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C8943 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# -0.00fF
C8944 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# 0.00fF
C8945 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# RESET_COUNTERn 0.02fF
C8946 sky130_fd_sc_hd__inv_1_35/Y RESET_COUNTERn 0.05fF
C8947 sky130_fd_sc_hd__dfrtn_1_28/a_761_289# sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C8948 sky130_fd_sc_hd__dfrtn_1_18/a_1270_413# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C8949 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C8950 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_2/a_805_47# 0.00fF
C8951 sky130_fd_sc_hd__dfrtn_1_42/a_761_289# sky130_fd_sc_hd__nor3_2_2/A 0.02fF
C8952 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_34/a_543_47# 0.00fF
C8953 sky130_fd_sc_hd__dfrtn_1_26/a_805_47# RESET_COUNTERn 0.00fF
C8954 sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C8955 sky130_fd_sc_hd__or2b_1_0/X sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C8956 sky130_fd_sc_hd__dfrtn_1_33/a_1217_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C8957 DOUT[9] sky130_fd_sc_hd__nor3_1_2/a_193_297# 0.00fF
C8958 VDD sky130_fd_sc_hd__inv_1_44/Y 0.53fF
C8959 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_3/a_639_47# 0.00fF
C8960 sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C8961 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# sky130_fd_sc_hd__dfrtp_1_3/a_1108_47# 0.00fF
C8962 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__dfrtp_1_3/a_651_413# 0.00fF
C8963 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__dfrtp_1_3/a_448_47# 0.00fF
C8964 sky130_fd_sc_hd__dfrtp_1_1/a_639_47# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C8965 sky130_fd_sc_hd__dfrtn_1_34/a_1217_47# RESET_COUNTERn -0.00fF
C8966 sky130_fd_sc_hd__dfrtn_1_16/a_639_47# sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C8967 sky130_fd_sc_hd__dfrtn_1_11/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C8968 sky130_fd_sc_hd__dfrtn_1_20/a_543_47# sky130_fd_sc_hd__dfrtn_1_21/a_1217_47# 0.00fF
C8969 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_21/a_761_289# 0.01fF
C8970 sky130_fd_sc_hd__dfrtn_1_20/a_761_289# sky130_fd_sc_hd__dfrtn_1_21/a_1270_413# 0.00fF
C8971 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__inv_1_43/A 0.45fF
C8972 sky130_fd_sc_hd__dfrtn_1_19/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_1108_47# -0.00fF
C8973 sky130_fd_sc_hd__dfrtn_1_36/a_543_47# sky130_fd_sc_hd__inv_1_40/A 0.00fF
C8974 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C8975 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C8976 sky130_fd_sc_hd__o2111a_2_0/X SEL_CONV_TIME[3] 0.03fF
C8977 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C8978 sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C8979 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_37/a_448_47# 0.00fF
C8980 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__dfrtn_1_37/a_193_47# 0.00fF
C8981 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_37/a_543_47# 0.00fF
C8982 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__dfrtn_1_37/a_761_289# 0.00fF
C8983 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_37/a_27_47# 0.00fF
C8984 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C8985 sky130_fd_sc_hd__mux4_2_0/X SEL_CONV_TIME[3] 0.02fF
C8986 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__nor3_2_0/A 0.01fF
C8987 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_2/a_543_47# 0.00fF
C8988 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C8989 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# 0.01fF
C8990 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_35/a_1270_413# 0.00fF
C8991 sky130_fd_sc_hd__inv_1_22/A sky130_fd_sc_hd__inv_1_23/A 0.24fF
C8992 sky130_fd_sc_hd__dfrtn_1_34/a_639_47# DONE 0.00fF
C8993 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__mux4_1_0/a_668_97# 0.00fF
C8994 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_24/a_761_289# -0.00fF
C8995 sky130_fd_sc_hd__nand2_1_0/a_113_47# DOUT[10] 0.00fF
C8996 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# 0.00fF
C8997 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# DOUT[2] 0.01fF
C8998 sky130_fd_sc_hd__nand2_1_2/a_113_47# SEL_CONV_TIME[1] 0.00fF
C8999 sky130_fd_sc_hd__dfrtn_1_27/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9000 DOUT[9] sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C9001 sky130_fd_sc_hd__dfrtn_1_38/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9002 sky130_fd_sc_hd__dfrtn_1_27/a_1217_47# VDD 0.00fF
C9003 sky130_fd_sc_hd__dfrtn_1_39/a_761_289# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C9004 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_18/a_1217_47# 0.00fF
C9005 DOUT[1] sky130_fd_sc_hd__dfrtn_1_22/a_1283_21# 0.00fF
C9006 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# DOUT[21] 0.00fF
C9007 SEL_CONV_TIME[2] sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C9008 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_41/a_27_47# 0.65fF
C9009 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# -0.00fF
C9010 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__nor3_1_0/a_193_297# 0.00fF
C9011 sky130_fd_sc_hd__dfrtn_1_26/a_761_289# DOUT[23] 0.00fF
C9012 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# DOUT[14] 0.00fF
C9013 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_3/a_193_47# 0.00fF
C9014 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__dfrtn_1_15/a_193_47# 0.00fF
C9015 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_543_47# 0.00fF
C9016 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_761_289# 0.00fF
C9017 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_15/a_27_47# 0.00fF
C9018 sky130_fd_sc_hd__mux4_2_0/X SEL_CONV_TIME[2] 0.02fF
C9019 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C9020 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C9021 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C9022 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C9023 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__inv_1_42/Y 0.27fF
C9024 sky130_fd_sc_hd__dfrtn_1_14/a_761_289# sky130_fd_sc_hd__nor3_1_0/a_109_297# 0.00fF
C9025 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__inv_1_54/Y 0.00fF
C9026 DOUT[16] sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C9027 sky130_fd_sc_hd__dfrtn_1_36/a_543_47# VDD 0.06fF
C9028 sky130_fd_sc_hd__dfrtn_1_36/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9029 sky130_fd_sc_hd__dfrtn_1_21/a_651_413# DOUT[2] 0.00fF
C9030 sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C9031 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# 0.00fF
C9032 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_543_47# 0.00fF
C9033 sky130_fd_sc_hd__dfrtn_1_0/a_651_413# DOUT[18] 0.00fF
C9034 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9035 sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9036 sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# sky130_fd_sc_hd__nor3_1_0/A 0.01fF
C9037 sky130_fd_sc_hd__dfrtn_1_17/a_543_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C9038 sky130_fd_sc_hd__dfrtn_1_12/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9039 sky130_fd_sc_hd__dfrtn_1_34/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9040 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_27/a_651_413# 0.00fF
C9041 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# 0.00fF
C9042 CLK_REF RESET_COUNTERn 0.34fF
C9043 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C9044 sky130_fd_sc_hd__dfrtn_1_28/a_1283_21# RESET_COUNTERn 0.01fF
C9045 sky130_fd_sc_hd__dfrtn_1_28/a_639_47# DOUT[21] 0.00fF
C9046 sky130_fd_sc_hd__dfrtn_1_14/a_651_413# sky130_fd_sc_hd__nor3_1_1/a_193_297# 0.00fF
C9047 sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C9048 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__or2_2_0/A 0.05fF
C9049 sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C9050 DOUT[4] sky130_fd_sc_hd__inv_1_48/A 0.01fF
C9051 sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# RESET_COUNTERn 0.00fF
C9052 sky130_fd_sc_hd__nor3_1_0/a_193_297# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C9053 sky130_fd_sc_hd__mux4_1_0/a_27_47# SEL_CONV_TIME[0] 0.00fF
C9054 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_11/a_761_289# 0.00fF
C9055 DOUT[1] sky130_fd_sc_hd__nor3_2_2/a_281_297# 0.00fF
C9056 sky130_fd_sc_hd__nor3_1_7/a_109_297# VDD 0.00fF
C9057 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C9058 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__inv_1_53/A 0.05fF
C9059 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__inv_1_4/Y 0.01fF
C9060 sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C9061 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_27_47# 0.00fF
C9062 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# SEL_CONV_TIME[2] 0.01fF
C9063 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C9064 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# VIN 0.00fF
C9065 sky130_fd_sc_hd__dfrtn_1_14/a_805_47# DOUT[22] 0.00fF
C9066 sky130_fd_sc_hd__inv_1_7/A DOUT[7] 0.00fF
C9067 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__inv_1_3/Y 0.02fF
C9068 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C9069 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C9070 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C9071 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C9072 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C9073 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C9074 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C9075 sky130_fd_sc_hd__dfrtn_1_40/a_1462_47# sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# 0.00fF
C9076 sky130_fd_sc_hd__dfrtn_1_32/a_543_47# sky130_fd_sc_hd__inv_1_9/A 0.01fF
C9077 sky130_fd_sc_hd__dfrtn_1_20/a_761_289# RESET_COUNTERn 0.01fF
C9078 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__inv_1_29/Y 0.21fF
C9079 sky130_fd_sc_hd__inv_1_4/A DOUT[19] 0.09fF
C9080 sky130_fd_sc_hd__dfrtn_1_18/a_543_47# DOUT[2] 0.01fF
C9081 DOUT[1] sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# 0.00fF
C9082 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C9083 sky130_fd_sc_hd__dfrtn_1_40/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9084 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__nor3_1_13/a_193_297# 0.00fF
C9085 sky130_fd_sc_hd__nor2_1_0/a_109_297# SEL_CONV_TIME[1] 0.00fF
C9086 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_25/a_1270_413# 0.00fF
C9087 sky130_fd_sc_hd__dfrtn_1_22/a_639_47# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C9088 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# -0.00fF
C9089 sky130_fd_sc_hd__nor3_1_4/A DOUT[3] 0.00fF
C9090 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C9091 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C9092 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__inv_1_48/A 0.03fF
C9093 sky130_fd_sc_hd__dfrtn_1_38/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C9094 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# 0.00fF
C9095 sky130_fd_sc_hd__or3b_2_0/a_472_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9096 sky130_fd_sc_hd__dfrtn_1_31/a_448_47# SEL_CONV_TIME[1] 0.00fF
C9097 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__nor3_1_4/A 0.20fF
C9098 sky130_fd_sc_hd__mux4_1_0/a_277_47# RESET_COUNTERn 0.01fF
C9099 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# RESET_COUNTERn 0.00fF
C9100 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# 0.00fF
C9101 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_19/a_1270_413# 0.00fF
C9102 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_12/A 0.00fF
C9103 sky130_fd_sc_hd__inv_1_33/A sky130_fd_sc_hd__inv_1_53/A 0.27fF
C9104 sky130_fd_sc_hd__or3b_2_0/a_472_297# sky130_fd_sc_hd__dfrtn_1_31/a_193_47# 0.00fF
C9105 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_543_47# 0.00fF
C9106 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_31/a_1283_21# 0.00fF
C9107 sky130_fd_sc_hd__or3b_2_0/a_388_297# sky130_fd_sc_hd__dfrtn_1_31/a_761_289# 0.00fF
C9108 sky130_fd_sc_hd__dfrtn_1_21/a_1217_47# sky130_fd_sc_hd__inv_1_35/A 0.00fF
C9109 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# DOUT[19] 0.00fF
C9110 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# 0.00fF
C9111 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C9112 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# 0.00fF
C9113 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# 0.00fF
C9114 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# 0.00fF
C9115 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C9116 sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C9117 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C9118 sky130_fd_sc_hd__dfrtn_1_17/a_651_413# VDD 0.01fF
C9119 sky130_fd_sc_hd__dfrtn_1_28/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C9120 sky130_fd_sc_hd__dfrtn_1_25/a_1462_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C9121 SLC_0/a_919_243# outb 0.01fF
C9122 sky130_fd_sc_hd__dfrtn_1_3/a_639_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C9123 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__inv_1_54/Y 0.00fF
C9124 sky130_fd_sc_hd__dfrtn_1_36/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9125 sky130_fd_sc_hd__dfrtn_1_14/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9126 sky130_fd_sc_hd__nor3_1_2/a_109_297# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C9127 sky130_fd_sc_hd__dfrtn_1_32/a_193_47# sky130_fd_sc_hd__dfrtn_1_32/a_761_289# -0.00fF
C9128 sky130_fd_sc_hd__dfrtn_1_32/a_27_47# sky130_fd_sc_hd__dfrtn_1_32/a_543_47# -0.00fF
C9129 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# 0.00fF
C9130 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__o2111a_2_0/a_566_47# 0.00fF
C9131 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_13/a_639_47# 0.00fF
C9132 sky130_fd_sc_hd__inv_1_15/A DOUT[3] 0.01fF
C9133 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C9134 sky130_fd_sc_hd__dfrtn_1_22/a_543_47# sky130_fd_sc_hd__inv_1_37/A 0.02fF
C9135 sky130_fd_sc_hd__dfrtn_1_3/a_651_413# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C9136 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C9137 DOUT[13] sky130_fd_sc_hd__inv_1_38/A 0.00fF
C9138 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C9139 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.01fF
C9140 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C9141 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C9142 sky130_fd_sc_hd__nor3_1_11/a_109_297# sky130_fd_sc_hd__dfrtn_1_7/a_27_47# 0.00fF
C9143 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_15/A 0.00fF
C9144 sky130_fd_sc_hd__o311a_1_0/a_585_47# SEL_CONV_TIME[0] 0.00fF
C9145 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfrtn_1_41/a_27_47# 0.02fF
C9146 sky130_fd_sc_hd__dfrtn_1_31/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9147 outb out 0.00fF
C9148 sky130_fd_sc_hd__dfrtn_1_31/a_1108_47# VDD 0.09fF
C9149 sky130_fd_sc_hd__mux4_2_0/a_872_316# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C9150 sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# sky130_fd_sc_hd__nor3_1_1/a_109_297# 0.00fF
C9151 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C9152 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C9153 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__inv_1_42/A 0.04fF
C9154 sky130_fd_sc_hd__mux4_2_0/a_600_345# SEL_CONV_TIME[0] 0.01fF
C9155 DOUT[5] sky130_fd_sc_hd__inv_1_15/A 0.03fF
C9156 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__inv_1_40/A 0.02fF
C9157 sky130_fd_sc_hd__dfrtn_1_0/a_1270_413# RESET_COUNTERn 0.00fF
C9158 sky130_fd_sc_hd__dfrtn_1_35/a_1283_21# RESET_COUNTERn 0.01fF
C9159 sky130_fd_sc_hd__dfrtn_1_35/a_639_47# DOUT[21] 0.00fF
C9160 sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C9161 sky130_fd_sc_hd__dfrtn_1_3/a_1462_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C9162 sky130_fd_sc_hd__nor3_1_11/a_193_297# sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# 0.00fF
C9163 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# sky130_fd_sc_hd__dfrtn_1_31/a_543_47# -0.00fF
C9164 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C9165 sky130_fd_sc_hd__dfrtn_1_23/a_805_47# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C9166 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C9167 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C9168 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# DOUT[3] 0.00fF
C9169 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# 0.00fF
C9170 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_39/a_1270_413# 0.00fF
C9171 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_1217_47# 0.00fF
C9172 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_805_47# 0.00fF
C9173 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# 0.00fF
C9174 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__inv_1_47/A 0.00fF
C9175 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# RESET_COUNTERn 0.00fF
C9176 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C9177 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_639_47# 0.00fF
C9178 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C9179 sky130_fd_sc_hd__dfrtn_1_4/a_543_47# sky130_fd_sc_hd__inv_1_5/A 0.01fF
C9180 sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C9181 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_19/a_651_413# 0.00fF
C9182 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_19/a_448_47# 0.00fF
C9183 sky130_fd_sc_hd__dfrtn_1_0/a_651_413# DOUT[22] 0.00fF
C9184 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__inv_1_31/A 0.00fF
C9185 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__nor3_2_3/C 0.08fF
C9186 sky130_fd_sc_hd__dfrtn_1_41/a_639_47# SEL_CONV_TIME[0] 0.00fF
C9187 sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C9188 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C9189 sky130_fd_sc_hd__dfrtn_1_34/a_543_47# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C9190 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_38/a_651_413# 0.00fF
C9191 sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# sky130_fd_sc_hd__inv_1_29/Y 0.00fF
C9192 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C9193 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_18/a_1270_413# 0.00fF
C9194 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# 0.00fF
C9195 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_805_47# 0.00fF
C9196 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C9197 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_1217_47# 0.00fF
C9198 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__dfrtn_1_18/a_761_289# 0.00fF
C9199 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C9200 sky130_fd_sc_hd__dfrtn_1_42/a_1270_413# sky130_fd_sc_hd__inv_1_25/A 0.00fF
C9201 sky130_fd_sc_hd__dfrtn_1_21/a_639_47# RESET_COUNTERn 0.00fF
C9202 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C9203 sky130_fd_sc_hd__dfrtn_1_32/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9204 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# 0.00fF
C9205 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# 0.00fF
C9206 sky130_fd_sc_hd__dfrtn_1_32/a_805_47# VDD 0.00fF
C9207 sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9208 sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C9209 sky130_fd_sc_hd__inv_1_13/A RESET_COUNTERn 0.18fF
C9210 sky130_fd_sc_hd__dfrtn_1_4/a_1270_413# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C9211 sky130_fd_sc_hd__or3_1_0/X sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C9212 sky130_fd_sc_hd__inv_1_42/A sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C9213 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_1/a_761_289# -0.00fF
C9214 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_1/a_543_47# -0.00fF
C9215 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# SEL_CONV_TIME[1] 0.02fF
C9216 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__nor3_1_19/Y 0.02fF
C9217 sky130_fd_sc_hd__dfrtn_1_36/a_1270_413# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C9218 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C9219 sky130_fd_sc_hd__o311a_1_0/a_266_47# DOUT[21] 0.00fF
C9220 sky130_fd_sc_hd__or3_1_0/a_183_297# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C9221 sky130_fd_sc_hd__dfrtp_1_3/a_448_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C9222 sky130_fd_sc_hd__inv_1_6/Y DOUT[7] 0.85fF
C9223 sky130_fd_sc_hd__dfrtn_1_27/a_761_289# SEL_CONV_TIME[0] 0.00fF
C9224 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9225 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C9226 sky130_fd_sc_hd__mux4_2_0/a_788_316# DOUT[21] 0.00fF
C9227 sky130_fd_sc_hd__or2b_1_0/a_301_297# VDD 0.00fF
C9228 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_26/a_639_47# 0.00fF
C9229 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C9230 VDD sky130_fd_sc_hd__inv_1_52/Y 0.76fF
C9231 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_24/a_639_47# 0.00fF
C9232 sky130_fd_sc_hd__dfrtn_1_25/a_1270_413# sky130_fd_sc_hd__dfrtn_1_28/a_27_47# 0.00fF
C9233 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_36/a_543_47# 0.01fF
C9234 sky130_fd_sc_hd__nor3_1_15/a_193_297# DOUT[16] 0.00fF
C9235 sky130_fd_sc_hd__dfrtn_1_21/a_543_47# sky130_fd_sc_hd__dfrtn_1_19/a_1283_21# 0.00fF
C9236 sky130_fd_sc_hd__nor3_1_4/A DOUT[20] -0.00fF
C9237 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__inv_1_8/A 0.65fF
C9238 sky130_fd_sc_hd__dfrtn_1_34/a_805_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C9239 sky130_fd_sc_hd__dfrtn_1_14/a_761_289# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C9240 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C9241 sky130_fd_sc_hd__dfrtn_1_42/a_448_47# sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C9242 sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# DOUT[11] 0.01fF
C9243 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__dfrtn_1_33/a_193_47# -0.17fF
C9244 sky130_fd_sc_hd__dfrtn_1_35/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9245 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C9246 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# DOUT[9] 0.00fF
C9247 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# VDD 0.00fF
C9248 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__inv_1_33/A 0.01fF
C9249 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# RESET_COUNTERn 0.02fF
C9250 sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# 0.00fF
C9251 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# 0.00fF
C9252 sky130_fd_sc_hd__inv_1_27/A SEL_CONV_TIME[1] 0.01fF
C9253 sky130_fd_sc_hd__o311a_1_0/a_266_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C9254 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# VDD -0.22fF
C9255 DOUT[4] sky130_fd_sc_hd__dfrtn_1_30/a_1270_413# 0.00fF
C9256 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__nor3_1_5/A 0.00fF
C9257 sky130_fd_sc_hd__inv_1_22/A DOUT[10] 0.01fF
C9258 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__dfrtn_1_30/a_805_47# -0.00fF
C9259 sky130_fd_sc_hd__nand3b_1_0/a_53_93# RESET_COUNTERn 0.00fF
C9260 sky130_fd_sc_hd__o221ai_1_0/a_213_123# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C9261 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C9262 sky130_fd_sc_hd__inv_1_13/Y sky130_fd_sc_hd__inv_1_6/A 0.00fF
C9263 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__inv_1_8/Y 0.43fF
C9264 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C9265 sky130_fd_sc_hd__dfrtn_1_19/a_1108_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C9266 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# 0.00fF
C9267 sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C9268 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.01fF
C9269 SLC_0/a_919_243# sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C9270 sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C9271 sky130_fd_sc_hd__dfrtn_1_28/a_1217_47# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C9272 sky130_fd_sc_hd__dfrtn_1_25/a_1270_413# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C9273 sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C9274 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__o211a_1_1/X 0.01fF
C9275 sky130_fd_sc_hd__inv_1_15/A DOUT[20] 0.00fF
C9276 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__nor3_2_3/C 0.20fF
C9277 sky130_fd_sc_hd__dfrtn_1_27/a_193_47# DOUT[21] 0.00fF
C9278 sky130_fd_sc_hd__dfrtn_1_19/a_1283_21# sky130_fd_sc_hd__inv_1_35/Y 0.00fF
C9279 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# 0.00fF
C9280 sky130_fd_sc_hd__dfrtn_1_3/a_761_289# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C9281 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__inv_1_12/A 0.01fF
C9282 sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# RESET_COUNTERn 0.00fF
C9283 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_25/a_193_47# 0.00fF
C9284 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__dfrtn_1_25/a_27_47# 0.00fF
C9285 sky130_fd_sc_hd__dfrtp_1_3/a_651_413# sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# 0.00fF
C9286 sky130_fd_sc_hd__dfrtp_1_3/a_639_47# sky130_fd_sc_hd__dfrtn_1_17/a_761_289# 0.00fF
C9287 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# 0.00fF
C9288 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_805_47# 0.00fF
C9289 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C9290 sky130_fd_sc_hd__dfrtn_1_12/a_651_413# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C9291 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C9292 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.00fF
C9293 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# -0.00fF
C9294 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtp_1_2/a_448_47# -0.00fF
C9295 sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C9296 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C9297 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C9298 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__inv_1_7/A 0.02fF
C9299 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__inv_1_11/Y 0.04fF
C9300 sky130_fd_sc_hd__inv_1_53/A sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C9301 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__dfrtn_1_29/a_639_47# 0.00fF
C9302 sky130_fd_sc_hd__dfrtn_1_4/a_651_413# sky130_fd_sc_hd__inv_1_7/A 0.01fF
C9303 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C9304 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# 0.00fF
C9305 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__dfrtn_1_24/a_27_47# 0.00fF
C9306 DOUT[9] DOUT[11] 0.05fF
C9307 sky130_fd_sc_hd__dfrtp_1_3/a_805_47# VDD 0.00fF
C9308 sky130_fd_sc_hd__dfrtp_1_3/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9309 sky130_fd_sc_hd__nor3_1_7/a_109_297# DOUT[3] 0.00fF
C9310 sky130_fd_sc_hd__inv_1_43/A RESET_COUNTERn 0.38fF
C9311 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__inv_1_53/A 0.01fF
C9312 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__inv_1_31/Y 0.01fF
C9313 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C9314 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.00fF
C9315 sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# SEL_CONV_TIME[1] 0.00fF
C9316 sky130_fd_sc_hd__nand3b_1_1/Y SEL_CONV_TIME[1] 0.16fF
C9317 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# VDD 0.10fF
C9318 sky130_fd_sc_hd__dfrtn_1_20/a_448_47# sky130_fd_sc_hd__dfrtn_1_21/a_193_47# 0.00fF
C9319 sky130_fd_sc_hd__dfrtn_1_21/a_651_413# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C9320 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C9321 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C9322 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__inv_1_43/Y 0.01fF
C9323 sky130_fd_sc_hd__nor3_2_3/a_27_297# sky130_fd_sc_hd__inv_1_39/Y 0.00fF
C9324 sky130_fd_sc_hd__inv_1_49/Y DOUT[13] 0.11fF
C9325 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__dfrtn_1_24/a_543_47# 0.00fF
C9326 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__dfrtn_1_24/a_761_289# 0.00fF
C9327 sky130_fd_sc_hd__dfrtn_1_28/a_543_47# sky130_fd_sc_hd__inv_1_48/A 0.01fF
C9328 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C9329 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C9330 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C9331 DOUT[4] sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# 0.01fF
C9332 sky130_fd_sc_hd__mux4_2_0/a_397_47# RESET_COUNTERn 0.00fF
C9333 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__inv_1_13/A 0.00fF
C9334 sky130_fd_sc_hd__dfrtp_1_1/a_448_47# sky130_fd_sc_hd__dfrtp_1_1/D -0.02fF
C9335 sky130_fd_sc_hd__dfrtn_1_23/a_761_289# sky130_fd_sc_hd__inv_1_40/A 0.01fF
C9336 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_651_413# -0.00fF
C9337 sky130_fd_sc_hd__dfrtn_1_11/a_639_47# RESET_COUNTERn 0.00fF
C9338 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_10/a_1283_21# 0.02fF
C9339 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# DOUT[23] 0.00fF
C9340 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# DOUT[19] 0.00fF
C9341 sky130_fd_sc_hd__dfrtn_1_8/a_1283_21# DOUT[12] 0.00fF
C9342 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_12/A 0.01fF
C9343 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__nor3_2_0/A 0.53fF
C9344 sky130_fd_sc_hd__nor3_1_0/a_193_297# DOUT[17] 0.00fF
C9345 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__or2b_1_0/X 0.01fF
C9346 sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# sky130_fd_sc_hd__inv_1_27/Y 0.00fF
C9347 sky130_fd_sc_hd__dfrtn_1_29/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9348 sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# VDD 0.00fF
C9349 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__inv_1_53/A 0.01fF
C9350 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_761_289# -0.00fF
C9351 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__dfrtp_1_3/a_543_47# -0.00fF
C9352 sky130_fd_sc_hd__dfrtp_1_2/a_805_47# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C9353 sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C9354 sky130_fd_sc_hd__dfrtp_1_1/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9355 DOUT[9] sky130_fd_sc_hd__nor3_1_5/a_109_297# 0.00fF
C9356 SEL_CONV_TIME[1] sky130_fd_sc_hd__inv_1_51/Y 0.01fF
C9357 CLK_REF sky130_fd_sc_hd__dfrtn_1_19/a_1283_21# 0.01fF
C9358 sky130_fd_sc_hd__dfrtp_1_2/a_639_47# sky130_fd_sc_hd__o211a_1_1/a_215_47# 0.00fF
C9359 sky130_fd_sc_hd__nor3_1_3/a_193_297# VDD 0.00fF
C9360 sky130_fd_sc_hd__dfrtn_1_20/a_805_47# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C9361 sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# sky130_fd_sc_hd__dfrtn_1_18/a_448_47# 0.00fF
C9362 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C9363 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__dfrtn_1_29/a_543_47# 0.00fF
C9364 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C9365 sky130_fd_sc_hd__dfrtn_1_18/a_543_47# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C9366 sky130_fd_sc_hd__nor3_1_16/a_193_297# sky130_fd_sc_hd__dfrtn_1_35/a_1283_21# 0.00fF
C9367 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C9368 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# DOUT[2] 0.01fF
C9369 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__nor3_2_1/A 0.12fF
C9370 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__o211a_1_0/a_510_47# 0.00fF
C9371 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# sky130_fd_sc_hd__o211a_1_0/a_79_21# 0.00fF
C9372 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# sky130_fd_sc_hd__dfrtn_1_36/a_448_47# 0.00fF
C9373 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__o211a_1_0/a_215_47# 0.00fF
C9374 sky130_fd_sc_hd__dfrtn_1_23/a_805_47# sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C9375 sky130_fd_sc_hd__dfrtn_1_23/a_639_47# sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C9376 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__inv_1_54/A 0.01fF
C9377 sky130_fd_sc_hd__dfrtn_1_27/a_651_413# RESET_COUNTERn 0.00fF
C9378 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_193_47# -0.03fF
C9379 sky130_fd_sc_hd__dfrtn_1_27/a_1462_47# DOUT[21] 0.00fF
C9380 sky130_fd_sc_hd__dfrtn_1_38/a_1270_413# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C9381 sky130_fd_sc_hd__or3b_2_0/X sky130_fd_sc_hd__inv_1_49/A 0.01fF
C9382 sky130_fd_sc_hd__dfrtn_1_35/a_1270_413# sky130_fd_sc_hd__inv_1_38/A 0.00fF
C9383 sky130_fd_sc_hd__nand3b_1_0/a_53_93# SEL_CONV_TIME[3] 0.02fF
C9384 sky130_fd_sc_hd__or2_2_0/a_39_297# DOUT[23] 0.00fF
C9385 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9386 sky130_fd_sc_hd__dfrtn_1_9/a_543_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C9387 sky130_fd_sc_hd__dfrtn_1_23/a_761_289# VDD 0.05fF
C9388 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__dfrtn_1_25/a_448_47# 0.00fF
C9389 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__dfrtn_1_25/a_805_47# 0.00fF
C9390 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_35/a_193_47# 0.00fF
C9391 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_32/a_805_47# 0.00fF
C9392 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C9393 sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C9394 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__dfrtn_1_34/a_543_47# -0.00fF
C9395 DOUT[13] DOUT[4] 0.23fF
C9396 DOUT[13] sky130_fd_sc_hd__dfrtn_1_30/a_543_47# 0.01fF
C9397 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C9398 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_761_289# 0.00fF
C9399 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C9400 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_543_47# 0.00fF
C9401 sky130_fd_sc_hd__dfrtn_1_38/a_448_47# DOUT[2] 0.00fF
C9402 sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.00fF
C9403 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# sky130_fd_sc_hd__mux4_2_0/a_1279_413# 0.00fF
C9404 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# sky130_fd_sc_hd__mux4_2_0/a_1060_369# 0.00fF
C9405 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# sky130_fd_sc_hd__mux4_2_0/a_397_47# 0.00fF
C9406 sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C9407 sky130_fd_sc_hd__mux4_2_0/a_1060_369# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9408 sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C9409 sky130_fd_sc_hd__dfrtn_1_10/a_1217_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C9410 sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# DOUT[21] 0.00fF
C9411 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# sky130_fd_sc_hd__inv_1_32/A 0.03fF
C9412 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# 0.00fF
C9413 DOUT[12] sky130_fd_sc_hd__inv_1_23/A 0.01fF
C9414 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__inv_1_8/A 0.00fF
C9415 DOUT[1] sky130_fd_sc_hd__inv_1_40/Y 0.22fF
C9416 sky130_fd_sc_hd__o221ai_1_0/a_109_47# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C9417 sky130_fd_sc_hd__inv_1_9/A DOUT[21] 0.01fF
C9418 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__or2_2_0/B 0.03fF
C9419 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# RESET_COUNTERn 0.00fF
C9420 sky130_fd_sc_hd__dfrtn_1_9/a_448_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C9421 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# 0.00fF
C9422 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# 0.00fF
C9423 DOUT[12] RESET_COUNTERn 0.01fF
C9424 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# sky130_fd_sc_hd__inv_1_0/Y 0.03fF
C9425 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# VDD 0.08fF
C9426 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9427 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C9428 sky130_fd_sc_hd__dfrtn_1_4/a_639_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C9429 sky130_fd_sc_hd__dfrtn_1_22/a_1462_47# VDD 0.00fF
C9430 sky130_fd_sc_hd__dfrtn_1_22/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9431 sky130_fd_sc_hd__nor3_1_12/a_193_297# sky130_fd_sc_hd__dfrtn_1_8/a_543_47# 0.00fF
C9432 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9433 sky130_fd_sc_hd__dfrtn_1_12/a_805_47# RESET_COUNTERn 0.00fF
C9434 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__nor3_1_1/a_193_297# 0.00fF
C9435 sky130_fd_sc_hd__dfrtn_1_38/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_651_413# -0.00fF
C9436 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_21/a_1462_47# 0.00fF
C9437 sky130_fd_sc_hd__dfrtn_1_20/a_805_47# sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# 0.00fF
C9438 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__inv_1_52/Y 0.02fF
C9439 DOUT[1] sky130_fd_sc_hd__dfrtn_1_42/a_805_47# 0.00fF
C9440 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C9441 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_33/A 0.00fF
C9442 VDD sky130_fd_sc_hd__inv_1_48/Y 0.23fF
C9443 sky130_fd_sc_hd__nand3b_1_0/a_232_47# sky130_fd_sc_hd__dfrtn_1_25/a_543_47# 0.00fF
C9444 sky130_fd_sc_hd__dfrtn_1_18/a_448_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C9445 sky130_fd_sc_hd__nor3_1_7/a_109_297# DOUT[20] 0.00fF
C9446 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C9447 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# 0.00fF
C9448 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/a_651_413# 0.00fF
C9449 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# sky130_fd_sc_hd__dfrtp_1_1/a_761_289# 0.00fF
C9450 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__mux4_2_0/a_1060_369# 0.00fF
C9451 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__mux4_2_0/a_872_316# 0.00fF
C9452 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.01fF
C9453 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C9454 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__dfrtn_1_13/a_27_47# 0.00fF
C9455 sky130_fd_sc_hd__dfrtn_1_26/a_448_47# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C9456 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_805_47# 0.00fF
C9457 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C9458 sky130_fd_sc_hd__mux4_2_0/a_397_47# SEL_CONV_TIME[3] 0.00fF
C9459 sky130_fd_sc_hd__dfrtn_1_3/a_1462_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C9460 sky130_fd_sc_hd__dfrtn_1_16/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9461 sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C9462 sky130_fd_sc_hd__dfrtn_1_16/a_805_47# VDD 0.00fF
C9463 sky130_fd_sc_hd__dfrtn_1_8/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C9464 sky130_fd_sc_hd__dfrtn_1_8/a_448_47# VDD 0.01fF
C9465 sky130_fd_sc_hd__nor3_1_18/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9466 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# -0.00fF
C9467 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# sky130_fd_sc_hd__dfrtn_1_29/a_543_47# -0.00fF
C9468 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# -0.00fF
C9469 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__inv_1_49/A 0.10fF
C9470 sky130_fd_sc_hd__dfrtn_1_7/a_651_413# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C9471 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C9472 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__inv_1_7/A 0.40fF
C9473 sky130_fd_sc_hd__a221oi_4_0/a_453_47# RESET_COUNTERn 0.00fF
C9474 sky130_fd_sc_hd__dfrtn_1_32/a_27_47# DOUT[21] 0.00fF
C9475 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_20/a_1270_413# 0.00fF
C9476 sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C9477 sky130_fd_sc_hd__inv_1_44/A sky130_fd_sc_hd__inv_1_48/A 0.00fF
C9478 DOUT[4] sky130_fd_sc_hd__dfrtn_1_10/a_27_47# 0.00fF
C9479 sky130_fd_sc_hd__dfrtn_1_31/a_651_413# SEL_CONV_TIME[0] 0.00fF
C9480 sky130_fd_sc_hd__nand3b_1_0/Y SEL_CONV_TIME[0] 0.42fF
C9481 sky130_fd_sc_hd__dfrtp_1_0/a_1462_47# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C9482 sky130_fd_sc_hd__inv_1_3/A RESET_COUNTERn 0.02fF
C9483 sky130_fd_sc_hd__nor3_1_12/a_109_297# RESET_COUNTERn 0.00fF
C9484 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C9485 sky130_fd_sc_hd__or3b_2_0/a_27_47# RESET_COUNTERn 0.03fF
C9486 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9487 sky130_fd_sc_hd__dfrtn_1_4/a_1270_413# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C9488 DOUT[1] sky130_fd_sc_hd__inv_1_36/Y 0.20fF
C9489 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# DOUT[14] 0.01fF
C9490 sky130_fd_sc_hd__dfrtn_1_9/a_651_413# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C9491 sky130_fd_sc_hd__mux4_2_0/a_397_47# SEL_CONV_TIME[2] 0.00fF
C9492 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# sky130_fd_sc_hd__or3_1_0/C 0.01fF
C9493 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# 0.00fF
C9494 sky130_fd_sc_hd__dfrtn_1_12/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9495 sky130_fd_sc_hd__o211a_1_1/a_215_47# sky130_fd_sc_hd__conb_1_0/LO 0.00fF
C9496 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.02fF
C9497 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# 0.00fF
C9498 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_38/a_1462_47# 0.00fF
C9499 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C9500 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_3/a_448_47# 0.00fF
C9501 sky130_fd_sc_hd__dfrtn_1_7/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9502 sky130_fd_sc_hd__dfrtn_1_7/a_639_47# VDD 0.00fF
C9503 sky130_fd_sc_hd__dfrtn_1_17/a_543_47# RESET_COUNTERn 0.01fF
C9504 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# sky130_fd_sc_hd__inv_1_54/A 0.01fF
C9505 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# DOUT[14] 0.00fF
C9506 sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C9507 sky130_fd_sc_hd__dfrtn_1_36/a_805_47# RESET_COUNTERn 0.00fF
C9508 sky130_fd_sc_hd__dfrtn_1_3/a_1270_413# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C9509 sky130_fd_sc_hd__dfrtn_1_21/a_639_47# sky130_fd_sc_hd__dfrtn_1_19/a_1283_21# 0.00fF
C9510 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_761_289# 0.00fF
C9511 DOUT[4] sky130_fd_sc_hd__dfrtn_1_28/a_1270_413# 0.00fF
C9512 sky130_fd_sc_hd__dfrtp_1_0/a_1462_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C9513 outb sky130_fd_sc_hd__inv_1_8/A 0.01fF
C9514 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__inv_1_7/A 0.02fF
C9515 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C9516 sky130_fd_sc_hd__dfrtn_1_11/a_761_289# sky130_fd_sc_hd__inv_1_11/Y 0.01fF
C9517 sky130_fd_sc_hd__nor3_2_3/C RESET_COUNTERn 2.83fF
C9518 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_543_47# 0.00fF
C9519 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C9520 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# 0.00fF
C9521 sky130_fd_sc_hd__mux4_2_0/a_1060_369# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C9522 VDD lc_out 5.28fF
C9523 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# RESET_COUNTERn 0.29fF
C9524 sky130_fd_sc_hd__dfrtn_1_20/a_761_289# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C9525 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C9526 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__nor3_1_4/A 0.01fF
C9527 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# sky130_fd_sc_hd__nor3_1_4/A 0.01fF
C9528 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C9529 sky130_fd_sc_hd__or2_2_0/a_121_297# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C9530 sky130_fd_sc_hd__or2_2_0/a_39_297# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C9531 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__inv_1_40/A 0.00fF
C9532 sky130_fd_sc_hd__dfrtn_1_27/a_805_47# DOUT[23] 0.00fF
C9533 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# 0.00fF
C9534 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C9535 sky130_fd_sc_hd__nor3_1_11/a_109_297# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C9536 sky130_fd_sc_hd__dfrtp_1_1/a_805_47# DOUT[0] 0.00fF
C9537 VDD DONE 1.70fF
C9538 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C9539 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C9540 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# SEL_CONV_TIME[1] 0.00fF
C9541 sky130_fd_sc_hd__dfrtn_1_25/a_651_413# sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# 0.00fF
C9542 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_805_47# 0.00fF
C9543 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# sky130_fd_sc_hd__dfrtn_1_27/a_1270_413# 0.00fF
C9544 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_1217_47# 0.00fF
C9545 sky130_fd_sc_hd__dfrtn_1_25/a_639_47# sky130_fd_sc_hd__dfrtn_1_27/a_761_289# 0.00fF
C9546 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_31/a_543_47# 0.00fF
C9547 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# DOUT[2] 0.01fF
C9548 sky130_fd_sc_hd__nor3_1_4/a_193_297# RESET_COUNTERn 0.00fF
C9549 sky130_fd_sc_hd__mux4_2_0/a_288_47# sky130_fd_sc_hd__inv_1_33/A 0.01fF
C9550 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C9551 sky130_fd_sc_hd__dfrtn_1_34/a_1462_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C9552 sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C9553 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C9554 sky130_fd_sc_hd__dfrtn_1_23/a_651_413# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C9555 sky130_fd_sc_hd__dfrtn_1_32/a_448_47# RESET_COUNTERn -0.00fF
C9556 sky130_fd_sc_hd__dfrtn_1_32/a_1217_47# DOUT[21] 0.00fF
C9557 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# SEL_CONV_TIME[0] 0.01fF
C9558 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__dfrtn_1_33/a_27_47# 0.00fF
C9559 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__dfrtn_1_33/a_543_47# 0.00fF
C9560 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_33/a_761_289# 0.00fF
C9561 sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__dfrtn_1_33/a_193_47# 0.00fF
C9562 sky130_fd_sc_hd__dfrtn_1_31/a_448_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C9563 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__dfrtn_1_14/a_543_47# -0.00fF
C9564 sky130_fd_sc_hd__dfrtn_1_8/a_1108_47# sky130_fd_sc_hd__inv_1_9/Y 0.00fF
C9565 sky130_fd_sc_hd__dfrtn_1_28/a_1283_21# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C9566 sky130_fd_sc_hd__dfrtp_1_2/a_805_47# CLK_REF 0.00fF
C9567 DOUT[4] sky130_fd_sc_hd__dfrtn_1_10/a_1217_47# 0.00fF
C9568 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__mux4_1_0/X 0.10fF
C9569 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C9570 sky130_fd_sc_hd__dfrtn_1_17/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9571 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# outb 0.00fF
C9572 sky130_fd_sc_hd__nor3_1_14/a_193_297# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C9573 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__dfrtn_1_22/a_651_413# -0.00fF
C9574 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# sky130_fd_sc_hd__dfrtn_1_22/a_448_47# -0.00fF
C9575 sky130_fd_sc_hd__dfrtn_1_36/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9576 sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C9577 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C9578 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C9579 sky130_fd_sc_hd__nand3b_1_1/a_232_47# SEL_CONV_TIME[1] 0.00fF
C9580 sky130_fd_sc_hd__a221oi_4_0/a_453_47# SEL_CONV_TIME[3] 0.01fF
C9581 sky130_fd_sc_hd__or3_1_0/a_111_297# SEL_CONV_TIME[1] 0.00fF
C9582 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__inv_1_14/A 0.01fF
C9583 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# VDD 0.08fF
C9584 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C9585 sky130_fd_sc_hd__inv_1_24/A outb 0.04fF
C9586 VDD sky130_fd_sc_hd__nor3_2_3/B 18.01fF
C9587 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_17/a_448_47# 0.00fF
C9588 sky130_fd_sc_hd__nor3_1_10/a_193_297# VDD 0.00fF
C9589 sky130_fd_sc_hd__dfrtn_1_39/a_639_47# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C9590 sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# VDD 0.10fF
C9591 sky130_fd_sc_hd__dfrtn_1_3/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C9592 sky130_fd_sc_hd__inv_1_7/A VIN 0.01fF
C9593 sky130_fd_sc_hd__dfrtn_1_14/a_761_289# sky130_fd_sc_hd__inv_1_1/A 0.01fF
C9594 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__inv_1_47/A 0.00fF
C9595 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_2/a_27_47# 0.00fF
C9596 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__inv_1_3/A 0.00fF
C9597 sky130_fd_sc_hd__nor3_1_3/a_193_297# DOUT[3] 0.00fF
C9598 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__or2b_1_0/a_219_297# 0.00fF
C9599 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__inv_1_47/A 0.01fF
C9600 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C9601 DOUT[9] sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C9602 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.01fF
C9603 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.01fF
C9604 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C9605 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C9606 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C9607 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# RESET_COUNTERn 0.01fF
C9608 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# sky130_fd_sc_hd__inv_1_51/Y 0.01fF
C9609 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C9610 sky130_fd_sc_hd__nand2_1_2/Y SEL_CONV_TIME[1] 0.06fF
C9611 sky130_fd_sc_hd__dfrtn_1_19/a_448_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C9612 sky130_fd_sc_hd__dfrtn_1_0/a_1462_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C9613 DOUT[4] sky130_fd_sc_hd__dfrtn_1_35/a_1270_413# 0.00fF
C9614 sky130_fd_sc_hd__nor3_1_3/a_193_297# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C9615 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# DOUT[21] 0.01fF
C9616 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# 0.00fF
C9617 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# 0.00fF
C9618 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_31/a_1283_21# 0.00fF
C9619 sky130_fd_sc_hd__a221oi_4_0/a_453_47# SEL_CONV_TIME[2] 0.01fF
C9620 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C9621 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C9622 sky130_fd_sc_hd__dfrtn_1_31/a_1462_47# RESET_COUNTERn 0.00fF
C9623 sky130_fd_sc_hd__nand3b_1_1/a_53_93# VDD 0.05fF
C9624 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# VDD -0.20fF
C9625 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_37/a_193_47# 0.00fF
C9626 sky130_fd_sc_hd__or3_1_0/a_29_53# VDD 0.07fF
C9627 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C9628 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__dfrtn_1_26/a_543_47# 0.01fF
C9629 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_26/a_761_289# 0.00fF
C9630 sky130_fd_sc_hd__o2111a_2_0/a_458_47# sky130_fd_sc_hd__dfrtn_1_28/a_27_47# 0.00fF
C9631 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_12/a_651_413# 0.00fF
C9632 sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C9633 sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9634 sky130_fd_sc_hd__dfrtn_1_25/a_651_413# SEL_CONV_TIME[1] 0.00fF
C9635 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C9636 sky130_fd_sc_hd__dfrtn_1_11/a_805_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C9637 sky130_fd_sc_hd__dfrtn_1_11/a_639_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C9638 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C9639 sky130_fd_sc_hd__nor3_2_3/C SEL_CONV_TIME[3] 0.22fF
C9640 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# 0.00fF
C9641 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__nor3_2_3/C 0.90fF
C9642 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_8/a_448_47# 0.00fF
C9643 sky130_fd_sc_hd__dfrtn_1_19/a_543_47# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C9644 sky130_fd_sc_hd__dfrtn_1_20/a_1217_47# DOUT[2] 0.00fF
C9645 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C9646 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# sky130_fd_sc_hd__dfrtn_1_16/a_543_47# -0.00fF
C9647 sky130_fd_sc_hd__dfrtn_1_16/a_193_47# sky130_fd_sc_hd__dfrtn_1_16/a_761_289# -0.00fF
C9648 sky130_fd_sc_hd__nor3_1_9/a_193_297# VDD 0.00fF
C9649 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# DOUT[3] 0.00fF
C9650 sky130_fd_sc_hd__dfrtn_1_31/a_805_47# DONE 0.00fF
C9651 sky130_fd_sc_hd__o221ai_1_0/a_213_123# sky130_fd_sc_hd__or2b_1_0/X 0.01fF
C9652 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C9653 sky130_fd_sc_hd__or2_2_0/B sky130_fd_sc_hd__o211a_1_1/X 0.00fF
C9654 sky130_fd_sc_hd__dfrtn_1_9/a_639_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C9655 sky130_fd_sc_hd__dfrtn_1_38/a_651_413# sky130_fd_sc_hd__inv_1_27/Y 0.00fF
C9656 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__o311a_1_0/A3 0.18fF
C9657 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__dfrtn_1_16/a_761_289# 0.00fF
C9658 sky130_fd_sc_hd__nor3_2_2/a_281_297# sky130_fd_sc_hd__dfrtn_1_16/a_193_47# 0.00fF
C9659 DOUT[12] DOUT[10] 0.04fF
C9660 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# sky130_fd_sc_hd__inv_1_2/A 0.02fF
C9661 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__dfrtn_1_33/a_1270_413# 0.00fF
C9662 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_33/a_805_47# 0.00fF
C9663 sky130_fd_sc_hd__nor3_1_19/Y sky130_fd_sc_hd__inv_1_42/A 0.00fF
C9664 sky130_fd_sc_hd__dfrtp_1_3/a_448_47# RESET_COUNTERn 0.00fF
C9665 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1_6/a_761_289# -0.00fF
C9666 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__o211a_1_1/a_215_47# 0.00fF
C9667 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__o211a_1_1/a_510_47# 0.00fF
C9668 sky130_fd_sc_hd__nor3_1_4/a_193_297# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C9669 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C9670 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__or2_2_0/B 0.01fF
C9671 sky130_fd_sc_hd__dfrtn_1_10/a_1217_47# outb 0.00fF
C9672 sky130_fd_sc_hd__or3_1_0/a_183_297# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C9673 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.02fF
C9674 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.02fF
C9675 sky130_fd_sc_hd__nor3_2_3/C SEL_CONV_TIME[2] 0.48fF
C9676 sky130_fd_sc_hd__o211a_1_0/X lc_out 0.00fF
C9677 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9678 sky130_fd_sc_hd__dfrtn_1_25/a_448_47# VDD 0.01fF
C9679 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C9680 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__dfrtn_1_3/a_193_47# 0.00fF
C9681 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__dfrtn_1_3/a_27_47# 0.01fF
C9682 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_3/a_761_289# 0.00fF
C9683 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__dfrtn_1_3/a_543_47# 0.00fF
C9684 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C9685 sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# sky130_fd_sc_hd__inv_1_35/Y 0.00fF
C9686 sky130_fd_sc_hd__nor3_1_4/a_109_297# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C9687 sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C9688 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C9689 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# DOUT[2] 0.01fF
C9690 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C9691 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__inv_1_13/A 0.00fF
C9692 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__or2_2_0/a_39_297# -0.00fF
C9693 sky130_fd_sc_hd__dfrtn_1_5/a_805_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C9694 sky130_fd_sc_hd__dfrtn_1_24/a_448_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C9695 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C9696 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# 0.00fF
C9697 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C9698 sky130_fd_sc_hd__nor3_1_15/a_193_297# RESET_COUNTERn 0.00fF
C9699 DOUT[1] sky130_fd_sc_hd__nor3_2_3/a_281_297# 0.00fF
C9700 sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# sky130_fd_sc_hd__inv_1_44/Y 0.02fF
C9701 VDD sky130_fd_sc_hd__nand2_1_1/Y 0.06fF
C9702 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__dfrtp_1_1/D 0.00fF
C9703 sky130_fd_sc_hd__dfrtn_1_42/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C9704 sky130_fd_sc_hd__nor3_1_7/a_193_297# DOUT[9] 0.00fF
C9705 sky130_fd_sc_hd__o211a_1_1/a_297_297# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C9706 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__or2_2_0/a_121_297# 0.00fF
C9707 sky130_fd_sc_hd__dfrtn_1_42/a_651_413# VDD 0.00fF
C9708 sky130_fd_sc_hd__o311a_1_0/a_266_297# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C9709 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C9710 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_7/A 0.00fF
C9711 sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# DOUT[21] 0.00fF
C9712 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# RESET_COUNTERn 0.00fF
C9713 sky130_fd_sc_hd__inv_1_37/A sky130_fd_sc_hd__inv_1_39/Y 0.12fF
C9714 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__inv_1_15/A 0.51fF
C9715 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C9716 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C9717 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C9718 DOUT[4] sky130_fd_sc_hd__inv_1_15/A 0.00fF
C9719 sky130_fd_sc_hd__nand3b_1_1/Y DOUT[21] 0.00fF
C9720 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C9721 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C9722 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_543_47# 0.00fF
C9723 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_761_289# 0.00fF
C9724 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C9725 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_36/a_651_413# 0.00fF
C9726 HEADER_0/a_508_138# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9727 sky130_fd_sc_hd__inv_1_6/Y VIN 0.10fF
C9728 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9729 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__o311a_1_0/a_266_297# 0.00fF
C9730 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# VDD 0.00fF
C9731 sky130_fd_sc_hd__nor3_1_3/a_193_297# DOUT[20] 0.00fF
C9732 sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C9733 sky130_fd_sc_hd__dfrtn_1_4/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9734 sky130_fd_sc_hd__dfrtn_1_38/a_639_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C9735 sky130_fd_sc_hd__dfrtn_1_14/a_639_47# DOUT[11] 0.00fF
C9736 sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# VDD 0.00fF
C9737 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_1/a_27_47# 0.00fF
C9738 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_1/a_193_47# 0.00fF
C9739 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# 0.00fF
C9740 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# 0.00fF
C9741 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_651_413# 0.00fF
C9742 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C9743 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.00fF
C9744 sky130_fd_sc_hd__or3b_2_0/a_388_297# sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C9745 sky130_fd_sc_hd__dfrtn_1_7/a_639_47# DOUT[3] 0.00fF
C9746 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C9747 SLC_0/a_264_22# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9748 SLC_0/a_1235_416# VDD 0.00fF
C9749 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# SEL_CONV_TIME[1] 0.00fF
C9750 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_193_47# -0.16fF
C9751 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C9752 sky130_fd_sc_hd__dfrtp_1_3/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9753 DOUT[23] sky130_fd_sc_hd__inv_1_38/Y 0.01fF
C9754 sky130_fd_sc_hd__o211a_1_0/X sky130_fd_sc_hd__nor3_2_3/B 0.13fF
C9755 sky130_fd_sc_hd__dfrtn_1_16/a_543_47# DOUT[15] 0.01fF
C9756 sky130_fd_sc_hd__dfrtn_1_33/a_761_289# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C9757 sky130_fd_sc_hd__dfrtn_1_7/a_639_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C9758 sky130_fd_sc_hd__dfrtn_1_8/a_27_47# sky130_fd_sc_hd__dfrtn_1_8/a_448_47# -0.00fF
C9759 sky130_fd_sc_hd__dfrtn_1_23/a_543_47# DOUT[21] 0.00fF
C9760 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__inv_1_45/Y 0.07fF
C9761 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C9762 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.00fF
C9763 sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C9764 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# sky130_fd_sc_hd__dfrtn_1_7/a_27_47# 0.00fF
C9765 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# 0.00fF
C9766 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# sky130_fd_sc_hd__dfrtn_1_7/a_543_47# 0.00fF
C9767 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_651_413# 0.00fF
C9768 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C9769 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# sky130_fd_sc_hd__nor3_1_4/a_193_297# 0.00fF
C9770 sky130_fd_sc_hd__nand3b_1_1/Y sky130_fd_sc_hd__o311a_1_0/A3 0.01fF
C9771 sky130_fd_sc_hd__inv_1_34/Y DOUT[2] 0.00fF
C9772 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__inv_1_0/Y 0.01fF
C9773 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_3/a_639_47# 0.00fF
C9774 DOUT[4] sky130_fd_sc_hd__dfrtn_1_12/a_543_47# 0.00fF
C9775 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_0/a_805_47# 0.00fF
C9776 sky130_fd_sc_hd__mux4_2_0/a_397_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C9777 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__dfrtn_1_28/a_1217_47# -0.00fF
C9778 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9779 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__inv_1_42/Y 0.01fF
C9780 sky130_fd_sc_hd__dfrtp_1_0/a_639_47# VDD 0.00fF
C9781 sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C9782 VDD DOUT[0] 3.25fF
C9783 sky130_fd_sc_hd__nor3_2_3/C DOUT[10] 0.03fF
C9784 sky130_fd_sc_hd__inv_1_51/Y DOUT[21] 0.00fF
C9785 sky130_fd_sc_hd__or3b_2_0/X sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C9786 sky130_fd_sc_hd__nand3b_1_0/a_232_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C9787 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# DOUT[7] 0.00fF
C9788 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# DOUT[6] 0.00fF
C9789 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# RESET_COUNTERn 0.15fF
C9790 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# DOUT[20] 0.00fF
C9791 sky130_fd_sc_hd__dfrtn_1_22/a_1270_413# RESET_COUNTERn 0.00fF
C9792 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.00fF
C9793 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_5/a_448_47# 0.00fF
C9794 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_639_47# 0.00fF
C9795 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C9796 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.00fF
C9797 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# 0.00fF
C9798 sky130_fd_sc_hd__dfrtn_1_39/a_805_47# VDD 0.00fF
C9799 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__nor3_2_3/B 0.20fF
C9800 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_32/a_543_47# 0.01fF
C9801 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__inv_1_44/A 0.01fF
C9802 sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9803 sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C9804 DOUT[4] sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C9805 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_10/a_448_47# -0.00fF
C9806 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# -0.00fF
C9807 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__dfrtn_1_3/a_639_47# 0.00fF
C9808 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# 0.00fF
C9809 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__dfrtn_1_3/a_1462_47# 0.00fF
C9810 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# 0.00fF
C9811 sky130_fd_sc_hd__dfrtn_1_11/a_761_289# outb 0.00fF
C9812 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9813 sky130_fd_sc_hd__dfrtn_1_18/a_805_47# VDD 0.00fF
C9814 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__dfrtn_1_25/a_639_47# 0.00fF
C9815 sky130_fd_sc_hd__inv_1_38/A sky130_fd_sc_hd__inv_1_52/Y 0.05fF
C9816 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C9817 sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# DOUT[2] 0.00fF
C9818 sky130_fd_sc_hd__o311a_1_0/A3 sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C9819 sky130_fd_sc_hd__dfrtn_1_17/a_193_47# sky130_fd_sc_hd__dfrtn_1_19/a_448_47# 0.00fF
C9820 sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# sky130_fd_sc_hd__dfrtn_1_19/a_543_47# 0.00fF
C9821 sky130_fd_sc_hd__dfrtn_1_17/a_651_413# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C9822 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# 0.00fF
C9823 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_43/A 0.00fF
C9824 sky130_fd_sc_hd__dfrtn_1_26/a_761_289# sky130_fd_sc_hd__inv_1_43/A 0.01fF
C9825 sky130_fd_sc_hd__dfrtn_1_16/a_448_47# RESET_COUNTERn 0.00fF
C9826 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# DOUT[14] 0.00fF
C9827 sky130_fd_sc_hd__or2_2_0/a_121_297# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C9828 sky130_fd_sc_hd__nor3_2_1/a_27_297# out 0.00fF
C9829 sky130_fd_sc_hd__dfrtn_1_8/a_761_289# RESET_COUNTERn 0.01fF
C9830 sky130_fd_sc_hd__dfrtn_1_8/a_651_413# DOUT[21] 0.00fF
C9831 sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9832 VDD sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.01fF
C9833 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_20/a_448_47# -0.00fF
C9834 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_20/a_651_413# -0.00fF
C9835 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__inv_1_30/Y 0.01fF
C9836 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# 0.00fF
C9837 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C9838 sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C9839 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# 0.00fF
C9840 sky130_fd_sc_hd__dfrtn_1_41/a_651_413# sky130_fd_sc_hd__dfrtn_1_38/a_651_413# 0.00fF
C9841 sky130_fd_sc_hd__dfrtn_1_32/a_193_47# sky130_fd_sc_hd__inv_1_36/Y 0.06fF
C9842 sky130_fd_sc_hd__nor3_1_14/a_193_297# DOUT[14] 0.00fF
C9843 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_13/a_27_47# 0.00fF
C9844 sky130_fd_sc_hd__dfrtn_1_19/a_448_47# VDD 0.01fF
C9845 sky130_fd_sc_hd__dfrtp_1_3/a_639_47# DOUT[23] 0.00fF
C9846 sky130_fd_sc_hd__nor3_2_3/B DOUT[3] 0.17fF
C9847 sky130_fd_sc_hd__nor3_1_10/a_193_297# DOUT[3] 0.00fF
C9848 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C9849 sky130_fd_sc_hd__nor3_1_13/a_109_297# sky130_fd_sc_hd__nor3_1_5/A 0.00fF
C9850 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__dfrtn_1_1/a_543_47# 0.00fF
C9851 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_1/a_639_47# 0.00fF
C9852 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C9853 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C9854 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_18/a_448_47# 0.00fF
C9855 sky130_fd_sc_hd__mux4_2_0/a_1064_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C9856 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__nor3_2_3/B 0.27fF
C9857 sky130_fd_sc_hd__nor3_1_10/a_193_297# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C9858 sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# SEL_CONV_TIME[1] 0.00fF
C9859 sky130_fd_sc_hd__dfrtn_1_31/a_543_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C9860 sky130_fd_sc_hd__dfrtn_1_31/a_448_47# sky130_fd_sc_hd__o221ai_1_0/a_295_297# 0.00fF
C9861 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_27/a_543_47# 0.00fF
C9862 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C9863 DOUT[4] sky130_fd_sc_hd__dfrtn_1_36/a_543_47# 0.00fF
C9864 DOUT[11] sky130_fd_sc_hd__inv_1_8/Y 0.01fF
C9865 DOUT[5] sky130_fd_sc_hd__nor3_2_3/B 0.03fF
C9866 sky130_fd_sc_hd__nor3_1_2/a_193_297# VDD 0.00fF
C9867 sky130_fd_sc_hd__dfrtp_1_2/a_639_47# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C9868 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C9869 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C9870 sky130_fd_sc_hd__dfrtn_1_23/a_639_47# RESET_COUNTERn 0.00fF
C9871 sky130_fd_sc_hd__dfrtn_1_22/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9872 sky130_fd_sc_hd__dfrtn_1_7/a_651_413# DOUT[7] 0.00fF
C9873 sky130_fd_sc_hd__dfrtn_1_7/a_639_47# DOUT[20] 0.00fF
C9874 sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# RESET_COUNTERn 0.00fF
C9875 sky130_fd_sc_hd__dfrtn_1_7/a_448_47# DOUT[8] 0.00fF
C9876 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# 0.00fF
C9877 sky130_fd_sc_hd__dfrtn_1_10/a_639_47# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C9878 sky130_fd_sc_hd__or3_1_0/X sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9879 sky130_fd_sc_hd__inv_1_31/Y SEL_CONV_TIME[1] 0.00fF
C9880 sky130_fd_sc_hd__inv_1_2/Y DOUT[14] 0.00fF
C9881 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# DOUT[3] 0.01fF
C9882 sky130_fd_sc_hd__dfrtn_1_30/a_761_289# sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.00fF
C9883 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# sky130_fd_sc_hd__dfrtn_1_0/a_651_413# -0.00fF
C9884 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# RESET_COUNTERn 0.00fF
C9885 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# DOUT[8] 0.00fF
C9886 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# CLK_REF 0.01fF
C9887 DOUT[7] RESET_COUNTERn 0.50fF
C9888 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C9889 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C9890 sky130_fd_sc_hd__dfrtn_1_14/a_761_289# DOUT[17] 0.00fF
C9891 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_1290_413# -0.01fF
C9892 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_750_97# -0.06fF
C9893 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C9894 sky130_fd_sc_hd__dfrtn_1_27/a_651_413# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C9895 sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.00fF
C9896 sky130_fd_sc_hd__dfrtn_1_26/a_639_47# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C9897 sky130_fd_sc_hd__nor3_1_9/a_193_297# DOUT[3] 0.00fF
C9898 HEADER_1/a_508_138# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C9899 sky130_fd_sc_hd__dfrtn_1_24/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9900 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__o311a_1_0/a_585_47# 0.00fF
C9901 sky130_fd_sc_hd__dfrtn_1_24/a_805_47# VDD 0.00fF
C9902 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C9903 sky130_fd_sc_hd__dfrtn_1_16/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C9904 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# VDD 0.05fF
C9905 sky130_fd_sc_hd__dfrtn_1_8/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C9906 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9907 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# sky130_fd_sc_hd__inv_1_36/A 0.01fF
C9908 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# SEL_CONV_TIME[0] 0.00fF
C9909 sky130_fd_sc_hd__inv_1_50/A RESET_COUNTERn 0.06fF
C9910 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C9911 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C9912 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C9913 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_31/a_1108_47# 0.00fF
C9914 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C9915 sky130_fd_sc_hd__dfrtn_1_9/a_639_47# DOUT[14] 0.00fF
C9916 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_12/a_193_47# 0.01fF
C9917 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__inv_1_14/A 0.05fF
C9918 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__mux4_2_0/a_872_316# 0.00fF
C9919 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_761_289# 0.00fF
C9920 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.02fF
C9921 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C9922 sky130_fd_sc_hd__o211a_1_1/a_215_47# sky130_fd_sc_hd__or2_2_0/A 0.01fF
C9923 CLK_REF sky130_fd_sc_hd__or2_2_0/a_39_297# 0.04fF
C9924 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_14/a_761_289# 0.00fF
C9925 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_14/a_193_47# 0.00fF
C9926 sky130_fd_sc_hd__dfrtn_1_30/a_805_47# SEL_CONV_TIME[1] 0.00fF
C9927 sky130_fd_sc_hd__dfrtn_1_20/a_1217_47# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C9928 sky130_fd_sc_hd__o211a_1_0/X DOUT[0] 0.01fF
C9929 sky130_fd_sc_hd__inv_1_12/A RESET_COUNTERn 0.30fF
C9930 sky130_fd_sc_hd__dfrtn_1_20/a_543_47# sky130_fd_sc_hd__dfrtn_1_21/a_27_47# 0.00fF
C9931 sky130_fd_sc_hd__dfrtn_1_23/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9932 sky130_fd_sc_hd__or3b_2_0/a_472_297# sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# 0.00fF
C9933 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_30/a_1270_413# 0.00fF
C9934 sky130_fd_sc_hd__inv_1_42/A SEL_CONV_TIME[0] 0.01fF
C9935 sky130_fd_sc_hd__nor3_2_2/A sky130_fd_sc_hd__nor3_2_3/C 1.04fF
C9936 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C9937 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# VDD 0.10fF
C9938 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__o221ai_1_0/a_493_297# 0.00fF
C9939 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_18/a_543_47# 0.00fF
C9940 sky130_fd_sc_hd__dfrtn_1_24/a_1462_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C9941 sky130_fd_sc_hd__dfrtn_1_7/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9942 sky130_fd_sc_hd__nand3b_1_1/a_316_47# SEL_CONV_TIME[0] 0.00fF
C9943 sky130_fd_sc_hd__or3_1_0/a_183_297# SEL_CONV_TIME[0] 0.00fF
C9944 sky130_fd_sc_hd__dfrtn_1_11/a_1270_413# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C9945 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C9946 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9947 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# VDD 0.06fF
C9948 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C9949 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C9950 sky130_fd_sc_hd__dfrtn_1_38/a_543_47# SEL_CONV_TIME[1] 0.00fF
C9951 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# RESET_COUNTERn -0.01fF
C9952 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C9953 sky130_fd_sc_hd__nor3_1_0/a_109_297# RESET_COUNTERn 0.00fF
C9954 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__dfrtn_1_30/a_761_289# 0.00fF
C9955 sky130_fd_sc_hd__nor3_2_3/B DOUT[20] 0.31fF
C9956 sky130_fd_sc_hd__nor3_1_10/a_109_297# DOUT[6] 0.00fF
C9957 sky130_fd_sc_hd__nor3_1_10/a_193_297# DOUT[20] 0.00fF
C9958 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_53/A 0.17fF
C9959 DOUT[15] sky130_fd_sc_hd__dfrtp_1_1/D 0.00fF
C9960 sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# VDD 0.10fF
C9961 sky130_fd_sc_hd__dfrtn_1_33/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C9962 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# RESET_COUNTERn 0.07fF
C9963 sky130_fd_sc_hd__dfrtn_1_22/a_543_47# sky130_fd_sc_hd__inv_1_40/Y 0.00fF
C9964 sky130_fd_sc_hd__dfrtn_1_30/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9965 sky130_fd_sc_hd__dfrtn_1_31/a_543_47# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C9966 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# DOUT[3] 0.00fF
C9967 sky130_fd_sc_hd__dfrtn_1_30/a_639_47# VDD 0.00fF
C9968 sky130_fd_sc_hd__inv_1_39/Y DOUT[14] 0.02fF
C9969 VDD DOUT[2] 2.98fF
C9970 sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# sky130_fd_sc_hd__inv_1_35/A 0.01fF
C9971 DOUT[4] sky130_fd_sc_hd__dfrtn_1_31/a_1108_47# 0.00fF
C9972 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C9973 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C9974 sky130_fd_sc_hd__dfrtn_1_30/a_651_413# sky130_fd_sc_hd__dfrtn_1_31/a_193_47# 0.00fF
C9975 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__dfrtn_1_31/a_651_413# 0.00fF
C9976 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__inv_1_11/A 0.01fF
C9977 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# DOUT[14] 0.00fF
C9978 sky130_fd_sc_hd__dfrtn_1_14/a_805_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C9979 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C9980 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_4/Y 0.01fF
C9981 sky130_fd_sc_hd__nor3_1_4/A sky130_fd_sc_hd__inv_1_13/Y 0.39fF
C9982 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# HEADER_0/a_508_138# 0.00fF
C9983 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__dfrtn_1_17/a_651_413# 0.00fF
C9984 sky130_fd_sc_hd__dfrtn_1_34/a_448_47# SEL_CONV_TIME[1] 0.00fF
C9985 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# 0.00fF
C9986 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C9987 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_29/a_543_47# 0.00fF
C9988 sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C9989 sky130_fd_sc_hd__nand3b_1_1/a_232_47# DOUT[21] 0.00fF
C9990 sky130_fd_sc_hd__or3_1_0/a_111_297# DOUT[21] 0.00fF
C9991 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C9992 sky130_fd_sc_hd__dfrtn_1_38/a_761_289# VDD 0.05fF
C9993 sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C9994 sky130_fd_sc_hd__nor3_2_0/A sky130_fd_sc_hd__inv_1_7/A 0.00fF
C9995 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__inv_1_45/A 0.36fF
C9996 sky130_fd_sc_hd__nor3_1_6/a_109_297# DOUT[9] 0.00fF
C9997 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# 0.01fF
C9998 sky130_fd_sc_hd__dfrtn_1_10/a_1283_21# sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# 0.00fF
C9999 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# 0.00fF
C10000 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# sky130_fd_sc_hd__dfrtn_1_11/a_193_47# 0.00fF
C10001 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_11/a_651_413# 0.00fF
C10002 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__dfrtn_1_11/a_761_289# 0.00fF
C10003 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_1270_413# 0.00fF
C10004 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C10005 sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C10006 sky130_fd_sc_hd__inv_1_7/Y DOUT[7] 0.00fF
C10007 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# DOUT[15] 0.00fF
C10008 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_12/a_1462_47# 0.00fF
C10009 DOUT[4] sky130_fd_sc_hd__dfrtn_1_32/a_805_47# 0.00fF
C10010 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# -0.00fF
C10011 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__dfrtp_1_1/a_543_47# -0.00fF
C10012 sky130_fd_sc_hd__dfrtn_1_12/a_639_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C10013 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__inv_1_40/Y 0.00fF
C10014 sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# sky130_fd_sc_hd__inv_1_6/A 0.01fF
C10015 sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# sky130_fd_sc_hd__dfrtn_1_17/a_761_289# 0.00fF
C10016 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_17/a_1270_413# 0.00fF
C10017 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# 0.00fF
C10018 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__dfrtn_1_17/a_805_47# 0.00fF
C10019 sky130_fd_sc_hd__dfrtp_1_2/a_805_47# sky130_fd_sc_hd__dfrtn_1_17/a_543_47# 0.00fF
C10020 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__dfrtn_1_40/a_1270_413# 0.00fF
C10021 sky130_fd_sc_hd__dfrtn_1_12/a_639_47# sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# 0.00fF
C10022 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# 0.00fF
C10023 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_4/Y 0.18fF
C10024 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__dfrtn_1_37/a_543_47# -0.00fF
C10025 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# -0.00fF
C10026 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C10027 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_14/a_651_413# 0.00fF
C10028 sky130_fd_sc_hd__dfrtn_1_28/a_1108_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C10029 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C10030 sky130_fd_sc_hd__dfrtn_1_26/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10031 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# VDD 0.08fF
C10032 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C10033 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# DOUT[14] 0.00fF
C10034 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__o2111a_2_0/a_80_21# 0.00fF
C10035 sky130_fd_sc_hd__or3_1_0/a_111_297# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C10036 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C10037 sky130_fd_sc_hd__inv_1_6/A DOUT[6] 0.01fF
C10038 sky130_fd_sc_hd__nor3_1_3/a_193_297# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C10039 sky130_fd_sc_hd__dfrtn_1_34/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10040 sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# VDD 0.08fF
C10041 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_7/a_761_289# 0.00fF
C10042 DOUT[4] sky130_fd_sc_hd__or2b_1_0/a_301_297# 0.00fF
C10043 sky130_fd_sc_hd__dfrtn_1_21/a_448_47# sky130_fd_sc_hd__dfrtn_1_21/a_27_47# -0.00fF
C10044 sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# VDD 0.00fF
C10045 sky130_fd_sc_hd__dfrtp_1_2/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10046 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# 0.00fF
C10047 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# 0.00fF
C10048 sky130_fd_sc_hd__inv_1_35/A sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C10049 sky130_fd_sc_hd__inv_1_24/A sky130_fd_sc_hd__inv_1_19/A 0.01fF
C10050 DOUT[4] sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C10051 sky130_fd_sc_hd__dfrtn_1_29/a_639_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C10052 sky130_fd_sc_hd__dfrtn_1_29/a_805_47# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C10053 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# sky130_fd_sc_hd__inv_1_40/Y 0.01fF
C10054 DOUT[9] sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C10055 sky130_fd_sc_hd__dfrtn_1_28/a_1108_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C10056 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_761_289# -0.00fF
C10057 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C10058 sky130_fd_sc_hd__o2111a_2_0/a_386_47# SEL_CONV_TIME[1] 0.00fF
C10059 sky130_fd_sc_hd__dfrtn_1_25/a_651_413# DOUT[21] 0.00fF
C10060 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# RESET_COUNTERn 0.01fF
C10061 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C10062 sky130_fd_sc_hd__dfrtp_1_1/a_639_47# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C10063 sky130_fd_sc_hd__dfrtn_1_37/a_1462_47# RESET_COUNTERn 0.00fF
C10064 sky130_fd_sc_hd__nor3_1_4/a_193_297# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C10065 sky130_fd_sc_hd__dfrtn_1_32/a_651_413# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C10066 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C10067 sky130_fd_sc_hd__nor3_1_19/a_193_297# SEL_CONV_TIME[1] 0.00fF
C10068 sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# RESET_COUNTERn 0.00fF
C10069 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__o311a_1_0/A3 0.01fF
C10070 sky130_fd_sc_hd__dfrtp_1_0/a_761_289# DOUT[15] 0.00fF
C10071 sky130_fd_sc_hd__or3b_2_0/a_388_297# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C10072 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.01fF
C10073 DOUT[4] sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C10074 DOUT[13] sky130_fd_sc_hd__or3b_2_0/a_176_21# 0.01fF
C10075 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__inv_1_43/A 0.01fF
C10076 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C10077 sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# HEADER_0/a_508_138# 0.00fF
C10078 sky130_fd_sc_hd__dfrtn_1_40/a_1270_413# VDD 0.00fF
C10079 sky130_fd_sc_hd__mux4_2_0/a_372_413# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C10080 sky130_fd_sc_hd__dfrtn_1_42/a_543_47# RESET_COUNTERn 0.02fF
C10081 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# SEL_CONV_TIME[3] 0.00fF
C10082 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C10083 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.00fF
C10084 sky130_fd_sc_hd__dfrtn_1_34/a_651_413# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C10085 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__inv_1_35/A 0.01fF
C10086 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C10087 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_10/a_543_47# 0.01fF
C10088 sky130_fd_sc_hd__dfrtn_1_0/a_651_413# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C10089 sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C10090 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C10091 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C10092 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__dfrtp_1_3/a_543_47# 0.00fF
C10093 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__mux4_2_0/a_193_369# -0.00fF
C10094 sky130_fd_sc_hd__dfrtp_1_1/a_639_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C10095 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# HEADER_0/a_508_138# 0.00fF
C10096 sky130_fd_sc_hd__dfrtn_1_0/a_805_47# DOUT[17] 0.00fF
C10097 sky130_fd_sc_hd__o2111a_2_0/a_674_297# VDD 0.00fF
C10098 HEADER_0/a_508_138# DOUT[7] 0.01fF
C10099 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# DOUT[7] 0.00fF
C10100 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# RESET_COUNTERn 0.02fF
C10101 sky130_fd_sc_hd__dfrtn_1_17/a_651_413# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C10102 sky130_fd_sc_hd__dfrtn_1_8/a_448_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C10103 sky130_fd_sc_hd__dfrtn_1_4/a_651_413# RESET_COUNTERn 0.00fF
C10104 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# SEL_CONV_TIME[0] 0.00fF
C10105 sky130_fd_sc_hd__dfrtn_1_33/a_1217_47# sky130_fd_sc_hd__inv_1_45/A 0.00fF
C10106 sky130_fd_sc_hd__inv_1_52/A DOUT[21] 0.00fF
C10107 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__dfrtn_1_34/a_193_47# 0.00fF
C10108 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__dfrtn_1_34/a_27_47# 0.00fF
C10109 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__nor3_1_3/a_109_297# 0.00fF
C10110 sky130_fd_sc_hd__nor3_1_19/a_109_297# VDD 0.00fF
C10111 sky130_fd_sc_hd__inv_1_26/A RESET_COUNTERn 0.25fF
C10112 sky130_fd_sc_hd__dfrtn_1_31/a_761_289# sky130_fd_sc_hd__inv_1_49/A 0.03fF
C10113 sky130_fd_sc_hd__dfrtn_1_42/a_1217_47# DOUT[15] 0.00fF
C10114 sky130_fd_sc_hd__nor3_1_2/a_193_297# DOUT[5] -0.00fF
C10115 DOUT[13] sky130_fd_sc_hd__dfrtn_1_31/a_27_47# 0.02fF
C10116 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# SEL_CONV_TIME[2] 0.02fF
C10117 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.26fF
C10118 sky130_fd_sc_hd__dfrtn_1_14/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C10119 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.05fF
C10120 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# VDD 0.07fF
C10121 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# 0.00fF
C10122 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C10123 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# 0.00fF
C10124 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# DOUT[3] 0.00fF
C10125 sky130_fd_sc_hd__dfrtp_1_0/a_1108_47# RESET_COUNTERn 0.02fF
C10126 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C10127 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__inv_1_45/Y 0.01fF
C10128 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_41/a_639_47# -0.00fF
C10129 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C10130 sky130_fd_sc_hd__o2111a_2_0/a_458_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C10131 sky130_fd_sc_hd__dfrtn_1_3/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10132 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_8/a_805_47# 0.00fF
C10133 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# lc_out 0.01fF
C10134 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C10135 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C10136 sky130_fd_sc_hd__dfrtn_1_39/a_448_47# RESET_COUNTERn 0.00fF
C10137 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C10138 sky130_fd_sc_hd__dfrtn_1_22/a_1283_21# sky130_fd_sc_hd__inv_1_39/Y 0.02fF
C10139 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__inv_1_13/A 0.61fF
C10140 sky130_fd_sc_hd__dfrtn_1_42/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.03fF
C10141 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# DOUT[21] 0.03fF
C10142 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__inv_1_8/Y 0.02fF
C10143 sky130_fd_sc_hd__dfrtp_1_3/a_639_47# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C10144 sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C10145 sky130_fd_sc_hd__inv_1_14/A RESET_COUNTERn 0.06fF
C10146 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__nor3_1_3/a_109_297# 0.00fF
C10147 sky130_fd_sc_hd__dfrtn_1_37/a_639_47# sky130_fd_sc_hd__inv_1_32/Y 0.00fF
C10148 DOUT[9] sky130_fd_sc_hd__nor3_1_1/a_109_297# 0.00fF
C10149 sky130_fd_sc_hd__dfrtn_1_18/a_448_47# RESET_COUNTERn 0.00fF
C10150 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__dfrtn_1_25/a_27_47# 0.00fF
C10151 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C10152 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# 0.00fF
C10153 sky130_fd_sc_hd__inv_1_38/A sky130_fd_sc_hd__nor3_2_3/B 0.08fF
C10154 en sky130_fd_sc_hd__inv_1_23/A 0.02fF
C10155 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10156 DOUT[4] sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# 0.00fF
C10157 sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10158 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# SEL_CONV_TIME[0] 0.05fF
C10159 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# SEL_CONV_TIME[3] 0.00fF
C10160 en RESET_COUNTERn 0.03fF
C10161 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_1270_413# 0.00fF
C10162 sky130_fd_sc_hd__inv_1_12/A DOUT[10] 0.01fF
C10163 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__nor3_2_0/a_281_297# 0.01fF
C10164 sky130_fd_sc_hd__dfrtn_1_37/a_1462_47# SEL_CONV_TIME[3] 0.00fF
C10165 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# DOUT[3] 0.00fF
C10166 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# VDD 0.09fF
C10167 sky130_fd_sc_hd__mux4_2_0/a_1064_47# sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.00fF
C10168 sky130_fd_sc_hd__mux4_2_0/a_872_316# sky130_fd_sc_hd__o311a_1_0/a_585_47# 0.00fF
C10169 sky130_fd_sc_hd__dfrtn_1_9/a_543_47# RESET_COUNTERn 0.01fF
C10170 VDD DOUT[11] 1.24fF
C10171 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__mux4_2_0/a_1060_369# -0.00fF
C10172 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C10173 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# 0.00fF
C10174 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# 0.00fF
C10175 sky130_fd_sc_hd__inv_1_44/Y sky130_fd_sc_hd__inv_1_44/A 0.38fF
C10176 sky130_fd_sc_hd__dfrtn_1_19/a_761_289# RESET_COUNTERn 0.02fF
C10177 CLK_REF sky130_fd_sc_hd__dfrtn_1_17/a_448_47# 0.00fF
C10178 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__inv_1_2/A 0.01fF
C10179 sky130_fd_sc_hd__mux4_2_0/a_372_413# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C10180 sky130_fd_sc_hd__dfrtn_1_24/a_1462_47# SEL_CONV_TIME[0] 0.00fF
C10181 sky130_fd_sc_hd__o221ai_1_0/a_213_123# RESET_COUNTERn 0.01fF
C10182 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__o2111a_2_0/a_566_47# 0.00fF
C10183 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10184 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_761_289# 0.00fF
C10185 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C10186 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C10187 sky130_fd_sc_hd__nor3_1_19/Y sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C10188 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__inv_1_8/A 0.02fF
C10189 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# -0.00fF
C10190 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C10191 sky130_fd_sc_hd__dfrtn_1_35/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# 0.00fF
C10192 sky130_fd_sc_hd__dfrtn_1_35/a_1108_47# DOUT[16] 0.00fF
C10193 sky130_fd_sc_hd__dfrtn_1_35/a_761_289# sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.00fF
C10194 sky130_fd_sc_hd__dfrtn_1_35/a_448_47# sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C10195 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# -0.00fF
C10196 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_25/a_448_47# -0.00fF
C10197 DOUT[13] sky130_fd_sc_hd__dfrtn_1_31/a_1217_47# 0.00fF
C10198 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_1270_413# 0.00fF
C10199 sky130_fd_sc_hd__dfrtn_1_37/a_1462_47# SEL_CONV_TIME[2] 0.00fF
C10200 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C10201 sky130_fd_sc_hd__dfrtn_1_28/a_639_47# VDD 0.00fF
C10202 sky130_fd_sc_hd__dfrtn_1_29/a_805_47# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C10203 sky130_fd_sc_hd__dfrtn_1_4/a_651_413# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C10204 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__inv_1_5/A 0.01fF
C10205 sky130_fd_sc_hd__dfrtn_1_25/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10206 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C10207 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# 0.02fF
C10208 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C10209 sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# sky130_fd_sc_hd__inv_1_12/A 0.02fF
C10210 sky130_fd_sc_hd__dfrtn_1_0/a_761_289# VDD 0.05fF
C10211 sky130_fd_sc_hd__dfrtn_1_7/a_1462_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C10212 sky130_fd_sc_hd__inv_1_9/Y sky130_fd_sc_hd__inv_1_8/A 0.26fF
C10213 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__nor3_2_3/B 0.31fF
C10214 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_1/Y 0.00fF
C10215 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__inv_1_48/A 0.01fF
C10216 sky130_fd_sc_hd__dfrtn_1_3/a_761_289# sky130_fd_sc_hd__inv_1_14/A 0.01fF
C10217 sky130_fd_sc_hd__mux4_1_0/a_27_47# SEL_CONV_TIME[1] 0.00fF
C10218 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_38/a_448_47# 0.00fF
C10219 VDD sky130_fd_sc_hd__nor3_1_5/a_109_297# 0.00fF
C10220 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C10221 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_14/a_193_47# 0.06fF
C10222 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__inv_1_6/A 0.01fF
C10223 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__nor3_2_3/C 0.35fF
C10224 sky130_fd_sc_hd__dfrtn_1_4/a_448_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C10225 sky130_fd_sc_hd__dfrtn_1_39/a_543_47# sky130_fd_sc_hd__inv_1_32/Y 0.00fF
C10226 sky130_fd_sc_hd__dfrtn_1_20/a_651_413# VDD 0.01fF
C10227 VDD sky130_fd_sc_hd__inv_1_30/Y 0.20fF
C10228 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C10229 sky130_fd_sc_hd__dfrtn_1_42/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10230 sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# DOUT[21] 0.00fF
C10231 sky130_fd_sc_hd__dfrtn_1_24/a_448_47# RESET_COUNTERn 0.00fF
C10232 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# RESET_COUNTERn 0.13fF
C10233 sky130_fd_sc_hd__dfrtn_1_25/a_639_47# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C10234 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C10235 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__nor3_2_3/B 0.34fF
C10236 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10237 sky130_fd_sc_hd__nor3_1_10/a_193_297# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C10238 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C10239 sky130_fd_sc_hd__dfrtn_1_20/a_805_47# sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# 0.00fF
C10240 DOUT[1] sky130_fd_sc_hd__dfrtn_1_36/a_651_413# 0.00fF
C10241 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C10242 sky130_fd_sc_hd__dfrtn_1_33/a_448_47# SEL_CONV_TIME[0] 0.00fF
C10243 sky130_fd_sc_hd__dfrtn_1_23/a_639_47# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C10244 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_12/a_193_47# -0.28fF
C10245 sky130_fd_sc_hd__dfrtn_1_16/a_1283_21# DOUT[2] 0.03fF
C10246 sky130_fd_sc_hd__dfrtn_1_42/a_193_47# sky130_fd_sc_hd__dfrtn_1_42/a_651_413# -0.00fF
C10247 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_193_47# 0.00fF
C10248 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_761_289# 0.00fF
C10249 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# sky130_fd_sc_hd__dfrtn_1_13/a_27_47# 0.00fF
C10250 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__inv_1_1/A 0.08fF
C10251 sky130_fd_sc_hd__o221ai_1_0/a_493_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10252 DOUT[9] sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C10253 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# DOUT[11] 0.00fF
C10254 sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# SEL_CONV_TIME[0] 0.00fF
C10255 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__dfrtp_1_0/a_193_47# -0.04fF
C10256 sky130_fd_sc_hd__inv_1_49/Y DONE 0.25fF
C10257 sky130_fd_sc_hd__mux4_1_0/a_1478_413# VDD 0.05fF
C10258 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C10259 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__inv_1_4/Y 0.01fF
C10260 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C10261 sky130_fd_sc_hd__dfrtn_1_10/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10262 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C10263 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C10264 sky130_fd_sc_hd__dfrtn_1_10/a_1462_47# VDD 0.00fF
C10265 sky130_fd_sc_hd__o211a_1_0/a_297_297# VDD 0.00fF
C10266 sky130_fd_sc_hd__dfrtn_1_11/a_761_289# sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# 0.00fF
C10267 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_639_47# 0.00fF
C10268 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# VIN 0.03fF
C10269 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__dfrtn_1_28/a_1283_21# 0.00fF
C10270 sky130_fd_sc_hd__dfrtp_1_0/a_1270_413# DOUT[23] 0.00fF
C10271 sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C10272 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_20/a_543_47# 0.00fF
C10273 DOUT[23] out 2.49fF
C10274 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_448_47# -0.00fF
C10275 sky130_fd_sc_hd__dfrtn_1_27/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# -0.00fF
C10276 sky130_fd_sc_hd__inv_1_54/A DOUT[23] 0.00fF
C10277 sky130_fd_sc_hd__nor3_1_15/a_109_297# DOUT[13] 0.00fF
C10278 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C10279 sky130_fd_sc_hd__inv_1_46/Y SEL_CONV_TIME[0] 0.00fF
C10280 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# 0.00fF
C10281 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C10282 sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C10283 sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# SEL_CONV_TIME[0] 0.00fF
C10284 sky130_fd_sc_hd__mux4_2_0/a_1279_413# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C10285 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_805_47# -0.00fF
C10286 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# DOUT[20] 0.00fF
C10287 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# DOUT[6] 0.00fF
C10288 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# RESET_COUNTERn 0.00fF
C10289 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_4/a_639_47# 0.00fF
C10290 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C10291 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# sky130_fd_sc_hd__dfrtn_1_4/a_543_47# 0.00fF
C10292 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__dfrtn_1_4/a_761_289# 0.00fF
C10293 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__dfrtn_1_4/a_448_47# 0.00fF
C10294 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_543_47# -0.00fF
C10295 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C10296 sky130_fd_sc_hd__dfrtn_1_39/a_448_47# SEL_CONV_TIME[2] 0.00fF
C10297 sky130_fd_sc_hd__inv_1_32/A sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C10298 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C10299 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.00fF
C10300 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__o311a_1_0/a_266_47# 0.00fF
C10301 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__o311a_1_0/a_368_297# 0.00fF
C10302 sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__inv_1_45/A 0.00fF
C10303 sky130_fd_sc_hd__or3b_2_0/X RESET_COUNTERn 0.11fF
C10304 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# RESET_COUNTERn 0.01fF
C10305 DOUT[1] sky130_fd_sc_hd__dfrtn_1_32/a_543_47# 0.00fF
C10306 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# DOUT[19] 0.00fF
C10307 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C10308 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C10309 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.00fF
C10310 sky130_fd_sc_hd__dfrtn_1_27/a_805_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C10311 sky130_fd_sc_hd__dfrtn_1_35/a_639_47# VDD 0.00fF
C10312 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__nor3_2_3/B 0.09fF
C10313 sky130_fd_sc_hd__dfrtn_1_12/a_639_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C10314 sky130_fd_sc_hd__o311a_1_0/a_585_47# SEL_CONV_TIME[1] 0.00fF
C10315 sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# RESET_COUNTERn 0.01fF
C10316 sky130_fd_sc_hd__dfrtn_1_21/a_761_289# sky130_fd_sc_hd__dfrtn_1_21/a_543_47# -0.00fF
C10317 sky130_fd_sc_hd__nor3_2_1/a_27_297# sky130_fd_sc_hd__o211a_1_0/a_79_21# 0.00fF
C10318 sky130_fd_sc_hd__inv_1_4/A DOUT[9] 0.02fF
C10319 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C10320 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.00fF
C10321 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C10322 SLC_0/a_264_22# sky130_fd_sc_hd__inv_1_26/A 0.00fF
C10323 sky130_fd_sc_hd__dfrtn_1_12/a_1462_47# DOUT[17] 0.00fF
C10324 sky130_fd_sc_hd__dfrtn_1_18/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_543_47# -0.00fF
C10325 sky130_fd_sc_hd__mux4_2_0/a_600_345# SEL_CONV_TIME[1] -0.00fF
C10326 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# DOUT[19] 0.00fF
C10327 sky130_fd_sc_hd__dfrtn_1_27/a_1270_413# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C10328 sky130_fd_sc_hd__dfrtn_1_34/a_651_413# SEL_CONV_TIME[0] 0.00fF
C10329 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__o221ai_1_0/a_295_297# 0.00fF
C10330 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10331 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# 0.00fF
C10332 sky130_fd_sc_hd__dfrtp_1_1/a_448_47# VDD 0.01fF
C10333 sky130_fd_sc_hd__dfrtn_1_23/a_805_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C10334 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_30/a_651_413# 0.00fF
C10335 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C10336 DOUT[4] DONE 0.03fF
C10337 sky130_fd_sc_hd__dfrtn_1_30/a_543_47# DONE 0.00fF
C10338 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C10339 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_805_47# -0.00fF
C10340 sky130_fd_sc_hd__dfrtp_1_0/a_1108_47# SLC_0/a_264_22# 0.00fF
C10341 sky130_fd_sc_hd__dfrtp_1_0/a_1283_21# SLC_0/a_919_243# 0.00fF
C10342 sky130_fd_sc_hd__dfrtn_1_16/a_193_47# sky130_fd_sc_hd__inv_1_25/A 0.00fF
C10343 sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# RESET_COUNTERn 0.00fF
C10344 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# sky130_fd_sc_hd__inv_1_26/A 0.00fF
C10345 sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10346 sky130_fd_sc_hd__nor3_1_17/a_193_297# DOUT[23] -0.00fF
C10347 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# DOUT[18] 0.00fF
C10348 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__nand3b_1_0/a_316_47# 0.00fF
C10349 CLK_REF sky130_fd_sc_hd__dfrtp_1_3/a_639_47# 0.00fF
C10350 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# 0.00fF
C10351 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# 0.00fF
C10352 sky130_fd_sc_hd__o211a_1_1/a_215_47# RESET_COUNTERn 0.00fF
C10353 sky130_fd_sc_hd__dfrtn_1_8/a_448_47# outb 0.00fF
C10354 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10355 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__inv_1_25/A 0.01fF
C10356 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_10/a_193_47# 0.24fF
C10357 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__dfrtn_1_13/a_651_413# 0.00fF
C10358 sky130_fd_sc_hd__o311a_1_0/a_266_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10359 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_12/a_448_47# 0.00fF
C10360 sky130_fd_sc_hd__dfrtn_1_7/a_651_413# VIN 0.01fF
C10361 sky130_fd_sc_hd__o311a_1_0/a_266_47# VDD 0.01fF
C10362 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfrtn_1_38/a_448_47# 0.00fF
C10363 sky130_fd_sc_hd__dfrtn_1_21/a_761_289# sky130_fd_sc_hd__inv_1_35/Y 0.01fF
C10364 DOUT[9] sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# 0.00fF
C10365 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C10366 sky130_fd_sc_hd__mux4_2_0/a_288_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C10367 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# DOUT[5] 0.00fF
C10368 sky130_fd_sc_hd__mux4_2_0/a_788_316# VDD 0.10fF
C10369 sky130_fd_sc_hd__dfrtp_1_0/a_1283_21# out 0.00fF
C10370 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C10371 sky130_fd_sc_hd__or2_2_0/a_39_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10372 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C10373 sky130_fd_sc_hd__inv_1_23/A VIN 0.85fF
C10374 sky130_fd_sc_hd__inv_1_4/Y DOUT[7] 0.46fF
C10375 sky130_fd_sc_hd__dfrtn_1_27/a_761_289# SEL_CONV_TIME[1] 0.00fF
C10376 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_2/a_27_47# 0.19fF
C10377 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# RESET_COUNTERn 0.08fF
C10378 sky130_fd_sc_hd__dfrtn_1_34/a_639_47# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C10379 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__inv_1_53/A 0.01fF
C10380 VIN RESET_COUNTERn 0.41fF
C10381 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# sky130_fd_sc_hd__inv_1_43/Y 0.07fF
C10382 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C10383 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__nand2_1_1/a_113_47# 0.00fF
C10384 sky130_fd_sc_hd__dfrtn_1_35/a_1283_21# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C10385 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10386 sky130_fd_sc_hd__o2111a_2_0/a_458_47# SEL_CONV_TIME[0] 0.00fF
C10387 sky130_fd_sc_hd__dfrtn_1_34/a_448_47# DOUT[21] 0.00fF
C10388 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# RESET_COUNTERn 0.01fF
C10389 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# VDD 0.05fF
C10390 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# RESET_COUNTERn 0.00fF
C10391 sky130_fd_sc_hd__dfrtn_1_35/a_543_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C10392 sky130_fd_sc_hd__nor3_1_20/a_193_297# VDD 0.00fF
C10393 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__nor3_2_3/B 0.31fF
C10394 DOUT[4] sky130_fd_sc_hd__nor3_2_3/B 0.20fF
C10395 sky130_fd_sc_hd__dfrtn_1_30/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10396 sky130_fd_sc_hd__dfrtn_1_41/a_1270_413# VDD 0.00fF
C10397 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C10398 sky130_fd_sc_hd__dfrtn_1_25/a_1462_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C10399 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# RESET_COUNTERn 0.00fF
C10400 sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# sky130_fd_sc_hd__inv_1_0/Y 0.01fF
C10401 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_34/a_543_47# 0.01fF
C10402 sky130_fd_sc_hd__dfrtn_1_8/a_193_47# sky130_fd_sc_hd__inv_1_8/A 0.13fF
C10403 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_39/a_639_47# 0.00fF
C10404 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__mux4_1_0/a_193_413# 0.00fF
C10405 DOUT[11] DOUT[3] 0.00fF
C10406 sky130_fd_sc_hd__nor3_1_11/a_109_297# DOUT[14] 0.00fF
C10407 sky130_fd_sc_hd__nor3_1_4/a_109_297# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C10408 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C10409 sky130_fd_sc_hd__dfrtn_1_33/a_1217_47# RESET_COUNTERn 0.00fF
C10410 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_30/a_1270_413# 0.00fF
C10411 en DOUT[10] 0.04fF
C10412 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# SEL_CONV_TIME[0] 0.00fF
C10413 sky130_fd_sc_hd__dfrtn_1_5/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10414 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C10415 sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C10416 sky130_fd_sc_hd__dfrtn_1_27/a_193_47# VDD 0.08fF
C10417 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# 0.00fF
C10418 sky130_fd_sc_hd__dfrtn_1_3/a_805_47# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.00fF
C10419 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# 0.00fF
C10420 sky130_fd_sc_hd__dfrtn_1_34/a_448_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C10421 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.29fF
C10422 sky130_fd_sc_hd__o211a_1_0/a_297_297# sky130_fd_sc_hd__o211a_1_0/X 0.00fF
C10423 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__dfrtn_1_1/a_27_47# 0.00fF
C10424 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# RESET_COUNTERn 0.01fF
C10425 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__inv_1_44/Y 0.01fF
C10426 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__inv_1_45/A 0.01fF
C10427 outb lc_out 0.00fF
C10428 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__inv_1_35/A 0.01fF
C10429 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10430 sky130_fd_sc_hd__dfrtn_1_17/a_1270_413# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C10431 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_193_47# -0.29fF
C10432 sky130_fd_sc_hd__dfrtn_1_37/a_639_47# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C10433 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C10434 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C10435 sky130_fd_sc_hd__o2111a_2_0/a_386_47# DOUT[21] 0.00fF
C10436 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C10437 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C10438 sky130_fd_sc_hd__o221ai_1_0/a_109_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C10439 sky130_fd_sc_hd__dfrtn_1_16/a_1462_47# sky130_fd_sc_hd__inv_1_25/A 0.00fF
C10440 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C10441 sky130_fd_sc_hd__or3b_2_0/a_388_297# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C10442 sky130_fd_sc_hd__dfrtn_1_38/a_639_47# RESET_COUNTERn 0.00fF
C10443 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__inv_1_43/Y 0.03fF
C10444 sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# DOUT[18] 0.00fF
C10445 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# 0.00fF
C10446 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_21/a_805_47# 0.00fF
C10447 CLK_REF sky130_fd_sc_hd__dfrtn_1_21/a_761_289# 0.00fF
C10448 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10449 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# VDD 0.03fF
C10450 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C10451 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C10452 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.00fF
C10453 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C10454 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_448_47# 0.00fF
C10455 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__inv_1_4/A 0.00fF
C10456 SEL_CONV_TIME[0] sky130_fd_sc_hd__mux4_1_0/X 0.06fF
C10457 sky130_fd_sc_hd__nor3_1_19/a_193_297# DOUT[21] 0.00fF
C10458 sky130_fd_sc_hd__dfrtp_1_3/a_543_47# sky130_fd_sc_hd__or2_2_0/B 0.02fF
C10459 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__inv_1_44/A 0.01fF
C10460 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# VDD 0.08fF
C10461 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_30/a_761_289# 0.00fF
C10462 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_10/a_1462_47# 0.00fF
C10463 sky130_fd_sc_hd__inv_1_0/A RESET_COUNTERn 0.34fF
C10464 sky130_fd_sc_hd__dfrtn_1_39/a_639_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C10465 sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# sky130_fd_sc_hd__inv_1_28/Y 0.01fF
C10466 sky130_fd_sc_hd__dfrtn_1_33/a_543_47# DOUT[23] 0.00fF
C10467 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10468 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__inv_1_19/A 0.04fF
C10469 sky130_fd_sc_hd__dfrtn_1_0/a_761_289# DOUT[5] 0.00fF
C10470 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# -0.00fF
C10471 sky130_fd_sc_hd__dfrtn_1_9/a_651_413# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C10472 VDD sky130_fd_sc_hd__inv_1_5/Y 0.39fF
C10473 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# RESET_COUNTERn -0.02fF
C10474 sky130_fd_sc_hd__dfrtn_1_28/a_543_47# sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C10475 sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# sky130_fd_sc_hd__dfrtn_1_13/a_27_47# 0.00fF
C10476 sky130_fd_sc_hd__dfrtn_1_42/a_543_47# sky130_fd_sc_hd__nor3_2_2/A 0.01fF
C10477 sky130_fd_sc_hd__o2111a_2_0/a_386_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C10478 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__inv_1_47/Y 0.00fF
C10479 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# 0.00fF
C10480 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# 0.01fF
C10481 sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# RESET_COUNTERn 0.00fF
C10482 sky130_fd_sc_hd__dfrtn_1_37/a_1462_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C10483 sky130_fd_sc_hd__dfrtn_1_33/a_1462_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C10484 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_639_47# 0.00fF
C10485 sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# sky130_fd_sc_hd__dfrtp_1_3/a_761_289# 0.00fF
C10486 sky130_fd_sc_hd__dfrtp_1_1/a_805_47# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C10487 sky130_fd_sc_hd__dfrtp_1_1/a_639_47# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C10488 sky130_fd_sc_hd__dfrtn_1_16/a_805_47# sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C10489 sky130_fd_sc_hd__inv_1_37/A DOUT[14] 0.71fF
C10490 sky130_fd_sc_hd__dfrtn_1_11/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10491 sky130_fd_sc_hd__dfrtn_1_34/a_1462_47# RESET_COUNTERn 0.00fF
C10492 sky130_fd_sc_hd__dfrtn_1_33/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10493 sky130_fd_sc_hd__dfrtn_1_20/a_543_47# sky130_fd_sc_hd__dfrtn_1_21/a_1270_413# 0.00fF
C10494 sky130_fd_sc_hd__nor3_1_5/a_109_297# DOUT[5] 0.00fF
C10495 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C10496 sky130_fd_sc_hd__dfrtn_1_19/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_448_47# -0.00fF
C10497 sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# sky130_fd_sc_hd__inv_1_40/A 0.00fF
C10498 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# DOUT[22] 0.00fF
C10499 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C10500 outb sky130_fd_sc_hd__nor3_2_3/B 0.35fF
C10501 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_37/a_193_47# 0.00fF
C10502 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_37/a_651_413# 0.00fF
C10503 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_37/a_27_47# 0.00fF
C10504 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__dfrtn_1_37/a_761_289# 0.00fF
C10505 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_37/a_448_47# 0.00fF
C10506 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C10507 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10508 sky130_fd_sc_hd__inv_1_1/A RESET_COUNTERn 0.47fF
C10509 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__nor3_2_0/A 0.01fF
C10510 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__dfrtn_1_2/a_543_47# 0.00fF
C10511 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# 0.00fF
C10512 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C10513 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_651_413# 0.00fF
C10514 sky130_fd_sc_hd__inv_1_7/Y VIN 0.01fF
C10515 sky130_fd_sc_hd__dfrtn_1_34/a_805_47# DONE 0.00fF
C10516 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__mux4_1_0/a_834_97# 0.00fF
C10517 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_24/a_761_289# -0.00fF
C10518 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_24/a_543_47# -0.00fF
C10519 sky130_fd_sc_hd__dfrtn_1_42/a_193_47# DOUT[2] 0.00fF
C10520 sky130_fd_sc_hd__inv_1_39/Y sky130_fd_sc_hd__inv_1_40/Y 0.01fF
C10521 sky130_fd_sc_hd__dfrtn_1_38/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10522 sky130_fd_sc_hd__dfrtn_1_27/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10523 sky130_fd_sc_hd__dfrtn_1_27/a_1462_47# VDD 0.00fF
C10524 sky130_fd_sc_hd__dfrtn_1_39/a_543_47# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C10525 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_18/a_1462_47# 0.00fF
C10526 DOUT[1] sky130_fd_sc_hd__dfrtn_1_22/a_1108_47# 0.00fF
C10527 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C10528 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_41/a_193_47# 0.59fF
C10529 sky130_fd_sc_hd__inv_1_28/A sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10530 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__nor3_2_0/A 0.01fF
C10531 sky130_fd_sc_hd__dfrtn_1_26/a_543_47# DOUT[23] 0.00fF
C10532 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# DOUT[14] 0.00fF
C10533 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_3/a_761_289# 0.00fF
C10534 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_543_47# 0.00fF
C10535 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__dfrtn_1_15/a_761_289# 0.00fF
C10536 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C10537 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_15/a_193_47# 0.00fF
C10538 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# sky130_fd_sc_hd__inv_1_42/Y 0.01fF
C10539 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C10540 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C10541 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_448_47# 0.00fF
C10542 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C10543 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C10544 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C10545 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__inv_1_54/Y 0.00fF
C10546 sky130_fd_sc_hd__dfrtn_1_14/a_761_289# sky130_fd_sc_hd__nor3_1_0/a_193_297# 0.00fF
C10547 sky130_fd_sc_hd__inv_1_1/Y DOUT[17] 0.00fF
C10548 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C10549 sky130_fd_sc_hd__dfrtn_1_36/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10550 DOUT[13] sky130_fd_sc_hd__or3b_2_0/B 0.01fF
C10551 sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# VDD 0.08fF
C10552 sky130_fd_sc_hd__dfrtn_1_21/a_193_47# DOUT[2] 0.00fF
C10553 sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C10554 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# 0.00fF
C10555 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# 0.00fF
C10556 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# SEL_CONV_TIME[3] 0.00fF
C10557 VDD sky130_fd_sc_hd__inv_1_9/A 1.04fF
C10558 sky130_fd_sc_hd__dfrtn_1_26/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10559 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10560 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C10561 sky130_fd_sc_hd__dfrtn_1_0/a_448_47# sky130_fd_sc_hd__nor3_1_0/A 0.01fF
C10562 sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C10563 sky130_fd_sc_hd__dfrtn_1_34/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10564 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C10565 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_1/a_639_47# 0.00fF
C10566 sky130_fd_sc_hd__nand2_1_2/a_113_47# VDD 0.00fF
C10567 sky130_fd_sc_hd__dfrtn_1_28/a_1108_47# RESET_COUNTERn 0.00fF
C10568 sky130_fd_sc_hd__dfrtn_1_28/a_805_47# DOUT[21] 0.00fF
C10569 sky130_fd_sc_hd__dfrtn_1_30/a_448_47# sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C10570 sky130_fd_sc_hd__dfrtn_1_39/a_448_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C10571 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# DOUT[9] 0.00fF
C10572 sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# RESET_COUNTERn 0.00fF
C10573 sky130_fd_sc_hd__mux4_1_0/a_193_47# SEL_CONV_TIME[0] 0.00fF
C10574 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_11/a_543_47# 0.00fF
C10575 sky130_fd_sc_hd__nor3_1_7/a_193_297# VDD 0.00fF
C10576 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_12/a_27_47# 0.00fF
C10577 sky130_fd_sc_hd__dfrtn_1_3/a_761_289# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C10578 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__inv_1_39/A 0.01fF
C10579 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C10580 HEADER_0/a_508_138# VIN 0.02fF
C10581 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_193_47# 0.00fF
C10582 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_27_47# 0.00fF
C10583 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# SEL_CONV_TIME[2] 0.05fF
C10584 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# VIN 0.00fF
C10585 sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.01fF
C10586 sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# DOUT[22] 0.00fF
C10587 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__inv_1_3/Y 0.02fF
C10588 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C10589 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_448_47# 0.00fF
C10590 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C10591 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C10592 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C10593 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C10594 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C10595 sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# sky130_fd_sc_hd__inv_1_9/A 0.00fF
C10596 sky130_fd_sc_hd__dfrtn_1_20/a_543_47# RESET_COUNTERn 0.01fF
C10597 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__inv_1_29/Y 0.01fF
C10598 DOUT[1] sky130_fd_sc_hd__dfrtn_1_23/a_448_47# 0.00fF
C10599 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.00fF
C10600 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C10601 sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# DOUT[2] 0.01fF
C10602 sky130_fd_sc_hd__dfrtn_1_32/a_27_47# VDD 0.20fF
C10603 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_25/a_639_47# 0.00fF
C10604 sky130_fd_sc_hd__inv_1_11/A RESET_COUNTERn 0.20fF
C10605 sky130_fd_sc_hd__dfrtn_1_22/a_805_47# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C10606 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# -0.00fF
C10607 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__inv_1_47/A 0.00fF
C10608 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C10609 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C10610 sky130_fd_sc_hd__o2111a_2_0/X sky130_fd_sc_hd__inv_1_48/A 0.00fF
C10611 sky130_fd_sc_hd__nor3_2_3/A sky130_fd_sc_hd__nor3_2_3/B 0.04fF
C10612 sky130_fd_sc_hd__dfrtn_1_31/a_651_413# SEL_CONV_TIME[1] 0.00fF
C10613 DOUT[1] DOUT[21] 0.02fF
C10614 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__inv_1_1/A 0.00fF
C10615 sky130_fd_sc_hd__nand3b_1_0/Y SEL_CONV_TIME[1] 0.02fF
C10616 sky130_fd_sc_hd__mux4_1_0/a_923_363# RESET_COUNTERn 0.00fF
C10617 VIN DOUT[10] 1.66fF
C10618 sky130_fd_sc_hd__dfrtn_1_10/a_1270_413# RESET_COUNTERn -0.00fF
C10619 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# 0.00fF
C10620 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__inv_1_48/A 0.00fF
C10621 HEADER_1/a_508_138# sky130_fd_sc_hd__inv_1_15/A 0.01fF
C10622 sky130_fd_sc_hd__or3b_2_0/a_388_297# sky130_fd_sc_hd__dfrtn_1_31/a_543_47# 0.00fF
C10623 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_1283_21# 0.00fF
C10624 sky130_fd_sc_hd__or3b_2_0/a_472_297# sky130_fd_sc_hd__dfrtn_1_31/a_761_289# 0.00fF
C10625 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_31/a_1108_47# 0.00fF
C10626 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_19/a_639_47# 0.00fF
C10627 sky130_fd_sc_hd__dfrtn_1_21/a_1270_413# sky130_fd_sc_hd__inv_1_35/A 0.00fF
C10628 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# DOUT[19] 0.00fF
C10629 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__inv_1_48/A 0.01fF
C10630 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# 0.00fF
C10631 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__dfrtn_1_15/a_639_47# 0.00fF
C10632 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C10633 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# 0.00fF
C10634 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# 0.00fF
C10635 sky130_fd_sc_hd__dfrtn_1_17/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10636 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# 0.00fF
C10637 sky130_fd_sc_hd__dfrtn_1_17/a_1270_413# VDD 0.00fF
C10638 sky130_fd_sc_hd__dfrtn_1_28/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.03fF
C10639 SLC_0/a_1235_416# outb 0.00fF
C10640 sky130_fd_sc_hd__dfrtn_1_3/a_805_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C10641 sky130_fd_sc_hd__dfrtn_1_14/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10642 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__nor3_1_0/a_109_297# 0.00fF
C10643 sky130_fd_sc_hd__nor2_1_0/a_109_297# VDD 0.00fF
C10644 sky130_fd_sc_hd__nor3_1_2/a_193_297# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C10645 sky130_fd_sc_hd__dfrtn_1_32/a_193_47# sky130_fd_sc_hd__dfrtn_1_32/a_543_47# -0.00fF
C10646 sky130_fd_sc_hd__nor3_2_3/a_281_297# sky130_fd_sc_hd__dfrtn_1_42/a_639_47# 0.00fF
C10647 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_13/a_805_47# 0.00fF
C10648 sky130_fd_sc_hd__dfrtn_1_22/a_1283_21# sky130_fd_sc_hd__inv_1_37/A 0.01fF
C10649 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__dfrtn_1_30/a_193_47# -0.03fF
C10650 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C10651 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C10652 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C10653 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.00fF
C10654 sky130_fd_sc_hd__nor3_1_11/a_109_297# sky130_fd_sc_hd__dfrtn_1_7/a_193_47# 0.00fF
C10655 sky130_fd_sc_hd__nor3_1_11/a_193_297# sky130_fd_sc_hd__dfrtn_1_7/a_27_47# 0.00fF
C10656 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfrtn_1_41/a_193_47# 0.22fF
C10657 sky130_fd_sc_hd__dfrtn_1_31/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10658 sky130_fd_sc_hd__dfrtn_1_31/a_448_47# VDD 0.01fF
C10659 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C10660 sky130_fd_sc_hd__mux4_2_0/a_1060_369# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C10661 sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# sky130_fd_sc_hd__nor3_1_1/a_193_297# 0.00fF
C10662 sky130_fd_sc_hd__dfrtn_1_38/a_193_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C10663 sky130_fd_sc_hd__dfrtn_1_28/a_193_47# sky130_fd_sc_hd__inv_1_42/A 0.28fF
C10664 sky130_fd_sc_hd__mux4_2_0/a_193_47# SEL_CONV_TIME[0] 0.00fF
C10665 sky130_fd_sc_hd__dfrtn_1_35/a_1108_47# RESET_COUNTERn 0.01fF
C10666 sky130_fd_sc_hd__dfrtn_1_35/a_805_47# DOUT[21] 0.00fF
C10667 sky130_fd_sc_hd__dfrtn_1_0/a_639_47# RESET_COUNTERn 0.00fF
C10668 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_1108_47# -0.00fF
C10669 sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C10670 sky130_fd_sc_hd__dfrtn_1_23/a_1217_47# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C10671 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C10672 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# DOUT[3] 0.00fF
C10673 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# 0.00fF
C10674 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_1462_47# 0.00fF
C10675 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_1217_47# 0.00fF
C10676 DOUT[19] sky130_fd_sc_hd__inv_1_2/Y 0.14fF
C10677 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_30/a_639_47# 0.00fF
C10678 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__inv_1_13/Y 0.14fF
C10679 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# RESET_COUNTERn 0.00fF
C10680 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C10681 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C10682 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_805_47# 0.00fF
C10683 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C10684 sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C10685 sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C10686 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__inv_1_31/A 0.00fF
C10687 sky130_fd_sc_hd__dfrtn_1_0/a_1270_413# DOUT[22] 0.00fF
C10688 sky130_fd_sc_hd__dfrtn_1_41/a_805_47# SEL_CONV_TIME[0] 0.00fF
C10689 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C10690 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_38/a_1270_413# 0.00fF
C10691 sky130_fd_sc_hd__dfrtn_1_34/a_543_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C10692 sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# sky130_fd_sc_hd__inv_1_29/Y 0.00fF
C10693 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C10694 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# 0.00fF
C10695 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_1217_47# 0.00fF
C10696 sky130_fd_sc_hd__dfrtn_1_40/a_1270_413# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C10697 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_1462_47# 0.00fF
C10698 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# sky130_fd_sc_hd__dfrtn_1_18/a_761_289# 0.00fF
C10699 sky130_fd_sc_hd__inv_1_50/Y sky130_fd_sc_hd__inv_1_49/A 0.01fF
C10700 sky130_fd_sc_hd__dfrtn_1_21/a_448_47# RESET_COUNTERn 0.01fF
C10701 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C10702 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.05fF
C10703 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C10704 sky130_fd_sc_hd__dfrtn_1_32/a_1217_47# VDD 0.00fF
C10705 sky130_fd_sc_hd__dfrtn_1_32/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10706 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C10707 sky130_fd_sc_hd__dfrtn_1_7/a_448_47# sky130_fd_sc_hd__inv_1_6/Y 0.01fF
C10708 sky130_fd_sc_hd__inv_1_5/Y DOUT[3] 0.02fF
C10709 sky130_fd_sc_hd__inv_1_39/A RESET_COUNTERn 0.12fF
C10710 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# VDD 0.14fF
C10711 sky130_fd_sc_hd__dfrtn_1_3/a_639_47# DOUT[11] 0.00fF
C10712 sky130_fd_sc_hd__dfrtn_1_4/a_639_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C10713 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_1/a_543_47# -0.00fF
C10714 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# -0.00fF
C10715 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# SEL_CONV_TIME[1] 0.00fF
C10716 sky130_fd_sc_hd__dfrtn_1_36/a_639_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C10717 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C10718 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_5/Y 0.03fF
C10719 sky130_fd_sc_hd__inv_1_6/Y DOUT[8] 0.24fF
C10720 sky130_fd_sc_hd__dfrtp_1_3/a_651_413# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C10721 sky130_fd_sc_hd__dfrtn_1_27/a_543_47# SEL_CONV_TIME[0] 0.00fF
C10722 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C10723 sky130_fd_sc_hd__mux4_2_0/a_27_47# RESET_COUNTERn 0.01fF
C10724 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10725 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_26/a_805_47# 0.00fF
C10726 sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C10727 sky130_fd_sc_hd__dfrtn_1_25/a_1270_413# sky130_fd_sc_hd__dfrtn_1_28/a_193_47# 0.00fF
C10728 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_24/a_805_47# 0.00fF
C10729 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.00fF
C10730 sky130_fd_sc_hd__nor3_1_15/a_193_297# sky130_fd_sc_hd__dfrtn_1_36/a_761_289# 0.00fF
C10731 sky130_fd_sc_hd__nor3_1_4/A DOUT[6] 0.00fF
C10732 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__inv_1_34/A 0.00fF
C10733 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__inv_1_9/A 0.01fF
C10734 sky130_fd_sc_hd__dfrtn_1_14/a_543_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C10735 sky130_fd_sc_hd__dfrtn_1_42/a_651_413# sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C10736 sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# DOUT[11] 0.01fF
C10737 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__dfrtn_1_33/a_761_289# -0.00fF
C10738 sky130_fd_sc_hd__dfrtn_1_0/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10739 sky130_fd_sc_hd__inv_1_35/A RESET_COUNTERn 0.12fF
C10740 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10741 sky130_fd_sc_hd__dfrtn_1_14/a_448_47# DOUT[9] 0.00fF
C10742 sky130_fd_sc_hd__dfrtn_1_35/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10743 sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# VDD 0.00fF
C10744 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__inv_1_33/A 0.01fF
C10745 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# RESET_COUNTERn 0.02fF
C10746 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# 0.00fF
C10747 DOUT[9] sky130_fd_sc_hd__inv_1_5/A 0.00fF
C10748 sky130_fd_sc_hd__o311a_1_0/a_585_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C10749 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# VDD 0.09fF
C10750 sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# sky130_fd_sc_hd__inv_1_15/A 0.01fF
C10751 DOUT[4] sky130_fd_sc_hd__dfrtn_1_30/a_639_47# 0.00fF
C10752 sky130_fd_sc_hd__nand3b_1_0/a_232_47# RESET_COUNTERn 0.00fF
C10753 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C10754 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C10755 DOUT[13] sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C10756 sky130_fd_sc_hd__dfrtn_1_19/a_448_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C10757 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# 0.00fF
C10758 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__o211a_1_1/a_297_297# 0.00fF
C10759 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.01fF
C10760 sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C10761 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C10762 sky130_fd_sc_hd__dfrtn_1_38/a_1462_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C10763 sky130_fd_sc_hd__dfrtn_1_28/a_1462_47# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C10764 sky130_fd_sc_hd__nor3_2_0/A RESET_COUNTERn 0.25fF
C10765 sky130_fd_sc_hd__dfrtn_1_25/a_639_47# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C10766 sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C10767 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__o211a_1_1/X 0.01fF
C10768 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.01fF
C10769 sky130_fd_sc_hd__dfrtn_1_27/a_761_289# DOUT[21] 0.00fF
C10770 sky130_fd_sc_hd__dfrtn_1_19/a_1108_47# sky130_fd_sc_hd__inv_1_35/Y 0.02fF
C10771 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# 0.00fF
C10772 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C10773 DOUT[17] RESET_COUNTERn 0.01fF
C10774 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C10775 sky130_fd_sc_hd__o211a_1_0/a_79_21# DOUT[23] 0.00fF
C10776 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_14/a_639_47# 0.00fF
C10777 sky130_fd_sc_hd__inv_1_44/A sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10778 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_25/a_761_289# 0.00fF
C10779 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__dfrtn_1_25/a_193_47# 0.00fF
C10780 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__dfrtn_1_25/a_27_47# 0.00fF
C10781 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_32/a_27_47# 0.00fF
C10782 sky130_fd_sc_hd__dfrtp_1_3/a_651_413# sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# 0.00fF
C10783 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_1462_47# 0.00fF
C10784 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# 0.00fF
C10785 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C10786 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtp_1_2/a_448_47# -0.00fF
C10787 sky130_fd_sc_hd__dfrtn_1_12/a_1270_413# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C10788 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.00fF
C10789 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C10790 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# sky130_fd_sc_hd__mux4_2_0/a_193_369# 0.00fF
C10791 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__mux4_2_0/a_372_413# 0.00fF
C10792 sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C10793 sky130_fd_sc_hd__inv_1_27/A VDD 1.05fF
C10794 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__inv_1_7/A 0.02fF
C10795 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C10796 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__inv_1_11/Y 0.09fF
C10797 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__dfrtn_1_29/a_639_47# 0.00fF
C10798 sky130_fd_sc_hd__dfrtn_1_4/a_1270_413# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C10799 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C10800 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# 0.00fF
C10801 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# sky130_fd_sc_hd__nor3_1_19/Y 0.01fF
C10802 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__dfrtn_1_24/a_193_47# 0.00fF
C10803 sky130_fd_sc_hd__or2_2_0/B sky130_fd_sc_hd__dfrtp_1_1/D 0.01fF
C10804 sky130_fd_sc_hd__dfrtp_1_3/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10805 sky130_fd_sc_hd__dfrtp_1_3/a_1217_47# VDD 0.00fF
C10806 sky130_fd_sc_hd__nor3_1_7/a_193_297# DOUT[3] 0.00fF
C10807 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__inv_1_31/Y 0.01fF
C10808 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.00fF
C10809 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_761_289# 0.00fF
C10810 sky130_fd_sc_hd__nor3_1_18/a_109_297# DOUT[15] 0.00fF
C10811 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10812 sky130_fd_sc_hd__dfrtn_1_22/a_761_289# VDD 0.05fF
C10813 DOUT[1] sky130_fd_sc_hd__dfrtn_1_42/a_27_47# 0.00fF
C10814 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# RESET_COUNTERn 0.06fF
C10815 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# 0.00fF
C10816 sky130_fd_sc_hd__dfrtn_1_20/a_651_413# sky130_fd_sc_hd__dfrtn_1_21/a_193_47# 0.00fF
C10817 sky130_fd_sc_hd__inv_1_45/Y sky130_fd_sc_hd__inv_1_43/Y 0.01fF
C10818 sky130_fd_sc_hd__dfrtn_1_21/a_193_47# sky130_fd_sc_hd__inv_1_30/Y 0.01fF
C10819 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__or2_2_0/a_121_297# 0.00fF
C10820 sky130_fd_sc_hd__nor3_2_3/a_281_297# sky130_fd_sc_hd__inv_1_39/Y 0.00fF
C10821 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__inv_1_43/Y 0.01fF
C10822 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__dfrtn_1_24/a_543_47# 0.00fF
C10823 sky130_fd_sc_hd__dfrtn_1_28/a_1283_21# sky130_fd_sc_hd__inv_1_48/A 0.01fF
C10824 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C10825 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C10826 DOUT[4] sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# 0.01fF
C10827 sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# 0.00fF
C10828 sky130_fd_sc_hd__mux4_2_0/a_1064_47# RESET_COUNTERn 0.00fF
C10829 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__inv_1_44/A 0.03fF
C10830 sky130_fd_sc_hd__nor3_1_3/a_109_297# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C10831 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C10832 sky130_fd_sc_hd__dfrtn_1_23/a_543_47# sky130_fd_sc_hd__inv_1_40/A 0.01fF
C10833 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C10834 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_639_47# -0.00fF
C10835 sky130_fd_sc_hd__inv_1_28/Y RESET_COUNTERn 0.03fF
C10836 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C10837 sky130_fd_sc_hd__dfrtn_1_11/a_805_47# RESET_COUNTERn 0.00fF
C10838 sky130_fd_sc_hd__dfrtn_1_8/a_27_47# sky130_fd_sc_hd__inv_1_9/A 0.00fF
C10839 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# 0.01fF
C10840 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C10841 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# DOUT[23] 0.00fF
C10842 sky130_fd_sc_hd__dfrtn_1_8/a_1108_47# DOUT[12] 0.00fF
C10843 sky130_fd_sc_hd__dfrtn_1_3/a_761_289# sky130_fd_sc_hd__nor3_2_0/A 0.02fF
C10844 sky130_fd_sc_hd__mux4_2_0/a_27_47# SEL_CONV_TIME[3] 0.02fF
C10845 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C10846 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# VDD -0.17fF
C10847 sky130_fd_sc_hd__inv_1_6/A sky130_fd_sc_hd__inv_1_13/A 0.00fF
C10848 sky130_fd_sc_hd__nor3_1_6/a_109_297# VDD 0.00fF
C10849 sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# sky130_fd_sc_hd__inv_1_27/Y 0.00fF
C10850 sky130_fd_sc_hd__dfrtn_1_29/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10851 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__inv_1_53/A 0.02fF
C10852 sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# VDD 0.00fF
C10853 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_543_47# -0.00fF
C10854 VDD sky130_fd_sc_hd__nand3b_1_1/Y 0.18fF
C10855 sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C10856 sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10857 DOUT[9] sky130_fd_sc_hd__nor3_1_5/a_193_297# 0.00fF
C10858 CLK_REF sky130_fd_sc_hd__dfrtn_1_19/a_1108_47# 0.01fF
C10859 sky130_fd_sc_hd__dfrtp_1_2/a_805_47# sky130_fd_sc_hd__o211a_1_1/a_215_47# 0.00fF
C10860 sky130_fd_sc_hd__nor3_1_3/a_109_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10861 sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# sky130_fd_sc_hd__dfrtn_1_18/a_651_413# 0.00fF
C10862 sky130_fd_sc_hd__dfrtn_1_20/a_1217_47# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C10863 sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# sky130_fd_sc_hd__dfrtn_1_18/a_448_47# 0.00fF
C10864 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C10865 sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C10866 sky130_fd_sc_hd__nor3_1_16/a_193_297# sky130_fd_sc_hd__dfrtn_1_35/a_1108_47# 0.00fF
C10867 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# DOUT[2] 0.00fF
C10868 sky130_fd_sc_hd__dfrtp_1_0/a_761_289# sky130_fd_sc_hd__nor3_2_1/A 0.01fF
C10869 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C10870 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# 0.00fF
C10871 sky130_fd_sc_hd__inv_1_4/Y VIN 0.04fF
C10872 sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# sky130_fd_sc_hd__dfrtn_1_36/a_448_47# 0.00fF
C10873 sky130_fd_sc_hd__dfrtn_1_23/a_1270_413# sky130_fd_sc_hd__dfrtn_1_36/a_543_47# 0.00fF
C10874 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__o211a_1_0/a_510_47# 0.00fF
C10875 sky130_fd_sc_hd__dfrtn_1_23/a_805_47# sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C10876 sky130_fd_sc_hd__dfrtn_1_23/a_1217_47# sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C10877 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# sky130_fd_sc_hd__dfrtn_1_36/a_651_413# 0.00fF
C10878 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__inv_1_54/A 0.01fF
C10879 sky130_fd_sc_hd__dfrtn_1_27/a_1270_413# RESET_COUNTERn 0.00fF
C10880 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_761_289# -0.00fF
C10881 sky130_fd_sc_hd__dfrtn_1_38/a_639_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C10882 CLK_REF sky130_fd_sc_hd__dfrtn_1_21/a_1462_47# 0.00fF
C10883 sky130_fd_sc_hd__dfrtn_1_35/a_639_47# sky130_fd_sc_hd__inv_1_38/A 0.00fF
C10884 sky130_fd_sc_hd__nand3b_1_0/a_232_47# SEL_CONV_TIME[3] 0.00fF
C10885 sky130_fd_sc_hd__or2_2_0/a_121_297# DOUT[23] 0.00fF
C10886 sky130_fd_sc_hd__mux4_2_0/a_27_47# SEL_CONV_TIME[2] 0.02fF
C10887 sky130_fd_sc_hd__nor3_1_11/a_109_297# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C10888 sky130_fd_sc_hd__dfrtn_1_23/a_543_47# VDD 0.06fF
C10889 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10890 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_35/a_761_289# 0.00fF
C10891 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_32/a_1217_47# 0.00fF
C10892 sky130_fd_sc_hd__nor3_2_3/C DOUT[18] 0.19fF
C10893 sky130_fd_sc_hd__dfrtn_1_30/a_448_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C10894 sky130_fd_sc_hd__nor3_2_0/a_27_297# sky130_fd_sc_hd__dfrtn_1_12/a_448_47# 0.00fF
C10895 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C10896 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# -0.00fF
C10897 sky130_fd_sc_hd__inv_1_43/Y sky130_fd_sc_hd__or3_1_0/C 0.00fF
C10898 DOUT[13] sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# 0.01fF
C10899 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C10900 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C10901 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_543_47# 0.00fF
C10902 sky130_fd_sc_hd__dfrtn_1_38/a_651_413# DOUT[2] 0.00fF
C10903 VDD sky130_fd_sc_hd__nor3_1_0/A 0.56fF
C10904 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__nor3_2_0/a_27_297# 0.01fF
C10905 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# sky130_fd_sc_hd__mux4_2_0/a_397_47# 0.00fF
C10906 sky130_fd_sc_hd__dfrtn_1_37/a_1462_47# sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.00fF
C10907 sky130_fd_sc_hd__dfrtn_1_42/a_1108_47# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C10908 sky130_fd_sc_hd__mux4_2_0/a_1279_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10909 sky130_fd_sc_hd__dfrtn_1_10/a_1462_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C10910 sky130_fd_sc_hd__dfrtn_1_22/a_1283_21# DOUT[14] 0.01fF
C10911 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# sky130_fd_sc_hd__inv_1_32/A 0.04fF
C10912 sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# DOUT[21] 0.00fF
C10913 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# RESET_COUNTERn 0.06fF
C10914 sky130_fd_sc_hd__nor3_1_19/Y SEL_CONV_TIME[0] 0.05fF
C10915 sky130_fd_sc_hd__o221ai_1_0/a_213_123# sky130_fd_sc_hd__inv_1_47/A 0.01fF
C10916 sky130_fd_sc_hd__inv_1_32/A sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10917 sky130_fd_sc_hd__inv_1_27/Y sky130_fd_sc_hd__inv_1_33/A 0.00fF
C10918 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# RESET_COUNTERn 0.00fF
C10919 sky130_fd_sc_hd__dfrtp_1_0/a_761_289# sky130_fd_sc_hd__or2_2_0/B 0.01fF
C10920 sky130_fd_sc_hd__dfrtn_1_9/a_651_413# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C10921 VDD sky130_fd_sc_hd__inv_1_51/Y 0.23fF
C10922 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# sky130_fd_sc_hd__inv_1_0/Y 0.01fF
C10923 sky130_fd_sc_hd__dfrtn_1_33/a_639_47# sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# 0.00fF
C10924 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# 0.00fF
C10925 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C10926 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# VDD 0.06fF
C10927 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# 0.00fF
C10928 sky130_fd_sc_hd__dfrtn_1_22/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10929 sky130_fd_sc_hd__dfrtn_1_39/a_651_413# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C10930 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_639_47# -0.00fF
C10931 DOUT[1] sky130_fd_sc_hd__dfrtn_1_42/a_1217_47# 0.00fF
C10932 sky130_fd_sc_hd__nor3_1_12/a_193_297# sky130_fd_sc_hd__dfrtn_1_8/a_1283_21# 0.00fF
C10933 sky130_fd_sc_hd__nor3_1_12/a_109_297# sky130_fd_sc_hd__dfrtn_1_8/a_1108_47# 0.00fF
C10934 sky130_fd_sc_hd__dfrtn_1_11/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10935 sky130_fd_sc_hd__dfrtn_1_12/a_1217_47# RESET_COUNTERn 0.00fF
C10936 sky130_fd_sc_hd__dfrtn_1_20/a_761_289# sky130_fd_sc_hd__dfrtn_1_21/a_1462_47# 0.00fF
C10937 sky130_fd_sc_hd__nor3_1_15/a_109_297# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C10938 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C10939 sky130_fd_sc_hd__nand3b_1_0/a_316_47# sky130_fd_sc_hd__dfrtn_1_25/a_543_47# 0.00fF
C10940 sky130_fd_sc_hd__dfrtn_1_26/a_639_47# DOUT[2] 0.00fF
C10941 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__inv_1_47/Y 0.00fF
C10942 sky130_fd_sc_hd__dfrtn_1_18/a_651_413# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C10943 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__o2111a_2_0/X 0.03fF
C10944 sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__inv_1_24/A 0.00fF
C10945 sky130_fd_sc_hd__nor3_1_7/a_193_297# DOUT[20] 0.00fF
C10946 sky130_fd_sc_hd__nor3_1_7/a_109_297# DOUT[6] 0.00fF
C10947 sky130_fd_sc_hd__inv_1_54/Y VDD 0.25fF
C10948 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C10949 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C10950 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# DOUT[23] 0.00fF
C10951 sky130_fd_sc_hd__dfrtp_1_0/a_639_47# sky130_fd_sc_hd__dfrtp_1_1/a_27_47# 0.00fF
C10952 sky130_fd_sc_hd__dfrtp_1_0/a_1108_47# sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# 0.00fF
C10953 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# sky130_fd_sc_hd__dfrtp_1_1/a_543_47# 0.00fF
C10954 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__dfrtp_1_1/a_639_47# 0.00fF
C10955 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# 0.00fF
C10956 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__mux4_2_0/a_872_316# 0.00fF
C10957 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__mux4_2_0/a_1279_413# 0.00fF
C10958 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# DOUT[0] 0.00fF
C10959 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C10960 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.01fF
C10961 sky130_fd_sc_hd__dfrtn_1_0/a_1217_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C10962 sky130_fd_sc_hd__dfrtn_1_8/a_1217_47# sky130_fd_sc_hd__inv_1_9/A 0.00fF
C10963 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C10964 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__dfrtn_1_13/a_193_47# 0.00fF
C10965 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__dfrtn_1_13/a_27_47# 0.00fF
C10966 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__inv_1_47/Y 0.00fF
C10967 sky130_fd_sc_hd__dfrtn_1_26/a_651_413# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C10968 sky130_fd_sc_hd__dfrtn_1_26/a_448_47# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C10969 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C10970 VDD DOUT[15] 10.82fF
C10971 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C10972 sky130_fd_sc_hd__mux4_2_0/a_1064_47# SEL_CONV_TIME[3] 0.00fF
C10973 sky130_fd_sc_hd__dfrtn_1_27/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C10974 sky130_fd_sc_hd__dfrtn_1_16/a_1217_47# VDD 0.00fF
C10975 sky130_fd_sc_hd__dfrtn_1_16/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C10976 sky130_fd_sc_hd__dfrtn_1_8/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C10977 sky130_fd_sc_hd__dfrtn_1_8/a_651_413# VDD 0.01fF
C10978 sky130_fd_sc_hd__nor3_1_18/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10979 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# sky130_fd_sc_hd__inv_1_49/A 0.02fF
C10980 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# -0.00fF
C10981 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_448_47# -0.00fF
C10982 sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C10983 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__inv_1_7/A 0.02fF
C10984 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# RESET_COUNTERn 0.00fF
C10985 DOUT[13] sky130_fd_sc_hd__dfrtn_1_34/a_27_47# 0.00fF
C10986 sky130_fd_sc_hd__dfrtn_1_24/a_448_47# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C10987 sky130_fd_sc_hd__dfrtn_1_32/a_193_47# DOUT[21] 0.00fF
C10988 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C10989 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# CLK_REF 0.02fF
C10990 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_20/a_639_47# 0.00fF
C10991 sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C10992 DOUT[4] sky130_fd_sc_hd__dfrtn_1_10/a_193_47# 0.00fF
C10993 sky130_fd_sc_hd__dfrtn_1_31/a_1270_413# SEL_CONV_TIME[0] 0.00fF
C10994 sky130_fd_sc_hd__nor3_1_12/a_193_297# RESET_COUNTERn 0.00fF
C10995 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C10996 sky130_fd_sc_hd__or3b_2_0/a_388_297# RESET_COUNTERn 0.00fF
C10997 sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C10998 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C10999 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# DOUT[14] 0.01fF
C11000 sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C11001 sky130_fd_sc_hd__mux4_2_0/a_1064_47# SEL_CONV_TIME[2] 0.00fF
C11002 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# sky130_fd_sc_hd__or3_1_0/C 0.01fF
C11003 sky130_fd_sc_hd__dfrtn_1_12/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11004 sky130_fd_sc_hd__or3_1_0/a_111_297# sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# 0.00fF
C11005 sky130_fd_sc_hd__or3_1_0/a_183_297# sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# 0.00fF
C11006 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__mux4_2_0/a_372_413# 0.00fF
C11007 sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C11008 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C11009 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_3/a_651_413# 0.00fF
C11010 sky130_fd_sc_hd__nor3_2_3/A DOUT[2] 0.03fF
C11011 sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11012 sky130_fd_sc_hd__dfrtn_1_7/a_805_47# VDD 0.00fF
C11013 sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# RESET_COUNTERn 0.05fF
C11014 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# sky130_fd_sc_hd__inv_1_54/A 0.01fF
C11015 sky130_fd_sc_hd__dfrtn_1_9/a_448_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C11016 sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# RESET_COUNTERn 0.00fF
C11017 sky130_fd_sc_hd__dfrtn_1_3/a_639_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C11018 sky130_fd_sc_hd__dfrtn_1_21/a_448_47# sky130_fd_sc_hd__dfrtn_1_19/a_1283_21# 0.00fF
C11019 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__inv_1_7/A 0.01fF
C11020 sky130_fd_sc_hd__dfrtn_1_0/a_761_289# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C11021 sky130_fd_sc_hd__nor3_1_1/a_109_297# VDD 0.00fF
C11022 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C11023 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# sky130_fd_sc_hd__inv_1_11/Y 0.02fF
C11024 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# 0.00fF
C11025 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_2/a_761_289# 0.00fF
C11026 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# 0.00fF
C11027 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C11028 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C11029 sky130_fd_sc_hd__dfrtn_1_31/a_761_289# RESET_COUNTERn 0.01fF
C11030 sky130_fd_sc_hd__nand3b_1_0/Y DOUT[21] 0.00fF
C11031 sky130_fd_sc_hd__dfrtn_1_20/a_543_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C11032 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__inv_1_13/Y 0.01fF
C11033 sky130_fd_sc_hd__dfrtn_1_9/a_761_289# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C11034 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11035 sky130_fd_sc_hd__or2_2_0/a_121_297# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C11036 sky130_fd_sc_hd__dfrtn_1_27/a_1217_47# DOUT[23] 0.00fF
C11037 DOUT[22] sky130_fd_sc_hd__nor3_2_3/C 0.75fF
C11038 sky130_fd_sc_hd__inv_1_37/A sky130_fd_sc_hd__inv_1_40/Y 0.02fF
C11039 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C11040 sky130_fd_sc_hd__nor3_1_11/a_193_297# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C11041 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C11042 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C11043 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# SEL_CONV_TIME[1] 0.00fF
C11044 sky130_fd_sc_hd__dfrtn_1_25/a_651_413# sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# 0.00fF
C11045 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_1462_47# 0.00fF
C11046 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_1217_47# 0.00fF
C11047 sky130_fd_sc_hd__dfrtn_1_25/a_1270_413# sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# 0.00fF
C11048 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# DOUT[2] 0.01fF
C11049 sky130_fd_sc_hd__o311a_1_0/a_368_297# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C11050 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# DONE 0.01fF
C11051 sky130_fd_sc_hd__nor3_1_10/a_109_297# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C11052 sky130_fd_sc_hd__mux4_2_0/a_372_413# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C11053 sky130_fd_sc_hd__dfrtn_1_19/a_1283_21# sky130_fd_sc_hd__inv_1_35/A 0.00fF
C11054 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11055 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__inv_1_43/A 0.01fF
C11056 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C11057 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C11058 DOUT[13] sky130_fd_sc_hd__dfrtn_1_34/a_1217_47# 0.00fF
C11059 sky130_fd_sc_hd__dfrtn_1_23/a_1270_413# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C11060 sky130_fd_sc_hd__dfrtn_1_32/a_651_413# RESET_COUNTERn 0.00fF
C11061 sky130_fd_sc_hd__dfrtn_1_32/a_1462_47# DOUT[21] 0.00fF
C11062 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# SEL_CONV_TIME[0] 0.01fF
C11063 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_33/a_543_47# 0.00fF
C11064 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__dfrtn_1_33/a_193_47# 0.00fF
C11065 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_33/a_27_47# 0.00fF
C11066 sky130_fd_sc_hd__dfrtn_1_31/a_651_413# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C11067 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__o311a_1_0/A3 0.12fF
C11068 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__nand2_1_1/a_113_47# 0.00fF
C11069 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# -0.00fF
C11070 sky130_fd_sc_hd__dfrtn_1_8/a_448_47# sky130_fd_sc_hd__inv_1_9/Y 0.01fF
C11071 sky130_fd_sc_hd__dfrtn_1_28/a_1108_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C11072 sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# CLK_REF 0.00fF
C11073 DOUT[4] sky130_fd_sc_hd__dfrtn_1_10/a_1462_47# 0.00fF
C11074 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__nand3b_1_1/a_53_93# 0.00fF
C11075 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__a221oi_4_0/a_471_297# 0.00fF
C11076 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# sky130_fd_sc_hd__inv_1_13/A 0.01fF
C11077 sky130_fd_sc_hd__dfrtn_1_17/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11078 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# sky130_fd_sc_hd__dfrtn_1_22/a_651_413# -0.00fF
C11079 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# outb 0.00fF
C11080 sky130_fd_sc_hd__inv_1_42/A SEL_CONV_TIME[1] 0.01fF
C11081 sky130_fd_sc_hd__dfrtn_1_36/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11082 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C11083 sky130_fd_sc_hd__dfrtn_1_24/a_805_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C11084 sky130_fd_sc_hd__nand3b_1_1/a_316_47# SEL_CONV_TIME[1] 0.00fF
C11085 sky130_fd_sc_hd__or3_1_0/a_183_297# SEL_CONV_TIME[1] 0.00fF
C11086 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# SEL_CONV_TIME[3] 0.01fF
C11087 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# VDD 0.01fF
C11088 sky130_fd_sc_hd__dfrtn_1_12/a_761_289# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C11089 sky130_fd_sc_hd__nor3_1_10/a_109_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11090 sky130_fd_sc_hd__nor3_1_6/a_109_297# DOUT[3] 0.00fF
C11091 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_17/a_651_413# 0.00fF
C11092 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C11093 sky130_fd_sc_hd__dfrtn_1_39/a_805_47# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C11094 sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# VDD 0.07fF
C11095 sky130_fd_sc_hd__dfrtn_1_14/a_543_47# sky130_fd_sc_hd__inv_1_1/A 0.01fF
C11096 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C11097 sky130_fd_sc_hd__nor3_1_16/a_109_297# DOUT[16] 0.00fF
C11098 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C11099 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_2/a_193_47# 0.00fF
C11100 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_2/a_27_47# 0.00fF
C11101 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__or2b_1_0/a_27_53# 0.00fF
C11102 DOUT[15] sky130_fd_sc_hd__o211a_1_0/X 0.07fF
C11103 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C11104 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__inv_1_47/A 0.02fF
C11105 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__nor3_1_4/A 0.01fF
C11106 sky130_fd_sc_hd__nand3b_1_0/a_232_47# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C11107 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# RESET_COUNTERn 0.01fF
C11108 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C11109 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C11110 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C11111 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C11112 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C11113 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C11114 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C11115 sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# sky130_fd_sc_hd__inv_1_38/A 0.00fF
C11116 sky130_fd_sc_hd__dfrtn_1_19/a_651_413# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C11117 DOUT[4] sky130_fd_sc_hd__dfrtn_1_35/a_639_47# 0.00fF
C11118 sky130_fd_sc_hd__nor3_2_2/A sky130_fd_sc_hd__inv_1_39/A 0.02fF
C11119 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# DOUT[21] 0.00fF
C11120 VDD sky130_fd_sc_hd__inv_1_32/Y 0.20fF
C11121 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_31/a_1108_47# 0.00fF
C11122 sky130_fd_sc_hd__nor3_1_4/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11123 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# SEL_CONV_TIME[2] 0.00fF
C11124 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C11125 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C11126 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__inv_1_43/Y 0.09fF
C11127 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_6/A 0.05fF
C11128 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_5/Y 0.01fF
C11129 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# sky130_fd_sc_hd__inv_1_5/Y 0.01fF
C11130 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# VDD 0.09fF
C11131 sky130_fd_sc_hd__nand3b_1_1/a_232_47# VDD 0.00fF
C11132 sky130_fd_sc_hd__or3_1_0/a_111_297# VDD 0.00fF
C11133 sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C11134 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# 0.00fF
C11135 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_26/a_543_47# 0.00fF
C11136 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__dfrtn_1_28/a_27_47# 0.00fF
C11137 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_12/a_1270_413# 0.00fF
C11138 sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11139 sky130_fd_sc_hd__nor3_2_1/a_27_297# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C11140 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C11141 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# 0.00fF
C11142 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_8/a_651_413# 0.00fF
C11143 sky130_fd_sc_hd__dfrtn_1_19/a_1283_21# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C11144 sky130_fd_sc_hd__dfrtn_1_20/a_1462_47# DOUT[2] 0.00fF
C11145 sky130_fd_sc_hd__dfrtn_1_16/a_193_47# sky130_fd_sc_hd__dfrtn_1_16/a_543_47# -0.00fF
C11146 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11147 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__dfrtn_1_23/a_639_47# 0.00fF
C11148 sky130_fd_sc_hd__dfrtn_1_22/a_639_47# sky130_fd_sc_hd__dfrtn_1_23/a_27_47# 0.00fF
C11149 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# DOUT[3] 0.00fF
C11150 sky130_fd_sc_hd__dfrtn_1_20/a_448_47# sky130_fd_sc_hd__dfrtn_1_21/a_543_47# 0.00fF
C11151 DOUT[5] sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C11152 sky130_fd_sc_hd__dfrtn_1_31/a_1217_47# DONE 0.00fF
C11153 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C11154 sky130_fd_sc_hd__dfrtn_1_9/a_805_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C11155 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# sky130_fd_sc_hd__o311a_1_0/A3 0.01fF
C11156 sky130_fd_sc_hd__dfrtn_1_38/a_1270_413# sky130_fd_sc_hd__inv_1_27/Y 0.00fF
C11157 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__nor3_1_4/A 0.01fF
C11158 sky130_fd_sc_hd__nand2_1_2/Y VDD 0.11fF
C11159 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_0/a_27_47# 0.65fF
C11160 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__inv_1_53/A 0.02fF
C11161 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__dfrtn_1_28/a_193_47# -0.15fF
C11162 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__dfrtn_1_16/a_543_47# 0.00fF
C11163 sky130_fd_sc_hd__nor3_2_2/a_281_297# sky130_fd_sc_hd__dfrtn_1_16/a_761_289# 0.00fF
C11164 DOUT[12] out 0.03fF
C11165 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__inv_1_2/A 0.02fF
C11166 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_33/a_1217_47# 0.00fF
C11167 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__dfrtn_1_33/a_448_47# 0.00fF
C11168 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_6/A 0.15fF
C11169 sky130_fd_sc_hd__inv_1_33/A sky130_fd_sc_hd__inv_1_44/Y 0.01fF
C11170 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C11171 sky130_fd_sc_hd__dfrtp_1_3/a_651_413# RESET_COUNTERn 0.00fF
C11172 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__dfrtn_1_6/a_761_289# -0.00fF
C11173 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1_6/a_543_47# -0.00fF
C11174 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C11175 sky130_fd_sc_hd__dfrtp_1_1/a_448_47# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.00fF
C11176 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__o211a_1_1/a_510_47# 0.00fF
C11177 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C11178 sky130_fd_sc_hd__dfrtn_1_10/a_1462_47# outb 0.00fF
C11179 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.00fF
C11180 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C11181 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C11182 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# VDD 0.27fF
C11183 sky130_fd_sc_hd__inv_1_35/A sky130_fd_sc_hd__inv_1_53/A 0.00fF
C11184 sky130_fd_sc_hd__inv_1_24/A sky130_fd_sc_hd__inv_1_22/A 0.01fF
C11185 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11186 sky130_fd_sc_hd__dfrtn_1_25/a_651_413# VDD 0.01fF
C11187 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C11188 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__dfrtn_1_3/a_27_47# 0.00fF
C11189 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__dfrtn_1_3/a_761_289# 0.00fF
C11190 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_3/a_543_47# 0.00fF
C11191 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__dfrtn_1_3/a_193_47# 0.00fF
C11192 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_448_47# 0.00fF
C11193 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C11194 sky130_fd_sc_hd__inv_1_4/A VDD 0.33fF
C11195 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_1_23/A 0.19fF
C11196 sky130_fd_sc_hd__dfrtn_1_18/a_27_47# VDD 0.20fF
C11197 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__inv_1_46/Y 0.00fF
C11198 sky130_fd_sc_hd__dfrtn_1_20/a_448_47# sky130_fd_sc_hd__inv_1_35/Y 0.00fF
C11199 sky130_fd_sc_hd__nor3_1_4/a_193_297# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C11200 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# DOUT[2] 0.00fF
C11201 sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# 0.00fF
C11202 sky130_fd_sc_hd__dfrtp_1_1/a_448_47# sky130_fd_sc_hd__dfrtp_1_2/a_448_47# 0.00fF
C11203 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__dfrtp_1_2/a_639_47# 0.00fF
C11204 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C11205 sky130_fd_sc_hd__inv_1_9/Y sky130_fd_sc_hd__nor3_2_3/B 0.06fF
C11206 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C11207 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_639_47# 0.00fF
C11208 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C11209 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C11210 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# sky130_fd_sc_hd__inv_1_44/Y 0.01fF
C11211 sky130_fd_sc_hd__o211a_1_1/a_215_47# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C11212 sky130_fd_sc_hd__dfrtn_1_42/a_1270_413# VDD 0.00fF
C11213 sky130_fd_sc_hd__dfrtn_1_42/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11214 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# DOUT[14] 0.02fF
C11215 sky130_fd_sc_hd__dfrtn_1_4/a_543_47# DOUT[14] 0.00fF
C11216 sky130_fd_sc_hd__o311a_1_0/a_368_297# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C11217 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_761_289# 0.00fF
C11218 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C11219 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C11220 sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# RESET_COUNTERn -0.00fF
C11221 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C11222 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C11223 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_543_47# 0.01fF
C11224 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# sky130_fd_sc_hd__dfrtn_1_38/a_761_289# 0.00fF
C11225 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.01fF
C11226 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__o311a_1_0/a_368_297# 0.00fF
C11227 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11228 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# VDD -0.00fF
C11229 sky130_fd_sc_hd__nor3_1_3/a_109_297# DOUT[7] 0.00fF
C11230 sky130_fd_sc_hd__dfrtn_1_4/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11231 sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C11232 sky130_fd_sc_hd__dfrtn_1_38/a_805_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C11233 sky130_fd_sc_hd__dfrtn_1_14/a_805_47# DOUT[11] 0.00fF
C11234 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_1/a_761_289# 0.00fF
C11235 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_1/a_193_47# 0.00fF
C11236 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_1/a_27_47# 0.00fF
C11237 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# 0.00fF
C11238 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# 0.00fF
C11239 sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__dfrtn_1_26/a_651_413# 0.00fF
C11240 sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# VDD 0.00fF
C11241 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__mux4_2_0/a_372_413# 0.00fF
C11242 sky130_fd_sc_hd__o311a_1_0/a_81_21# sky130_fd_sc_hd__inv_1_41/Y 0.04fF
C11243 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C11244 sky130_fd_sc_hd__or3b_2_0/a_472_297# sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C11245 sky130_fd_sc_hd__dfrtn_1_7/a_805_47# DOUT[3] 0.00fF
C11246 sky130_fd_sc_hd__inv_1_52/A VDD 1.44fF
C11247 sky130_fd_sc_hd__nor3_1_11/a_109_297# DOUT[19] 0.00fF
C11248 sky130_fd_sc_hd__dfrtn_1_19/a_543_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C11249 sky130_fd_sc_hd__nor3_1_14/a_109_297# VDD 0.00fF
C11250 SLC_0/a_919_243# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11251 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# SEL_CONV_TIME[1] 0.00fF
C11252 sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# VDD 0.10fF
C11253 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_761_289# -0.00fF
C11254 sky130_fd_sc_hd__dfrtp_1_3/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11255 sky130_fd_sc_hd__dfrtn_1_16/a_1283_21# DOUT[15] 0.01fF
C11256 sky130_fd_sc_hd__dfrtn_1_33/a_543_47# sky130_fd_sc_hd__inv_1_43/A 0.01fF
C11257 sky130_fd_sc_hd__dfrtn_1_7/a_805_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C11258 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# DOUT[21] 0.01fF
C11259 sky130_fd_sc_hd__dfrtn_1_8/a_27_47# sky130_fd_sc_hd__dfrtn_1_8/a_651_413# -0.00fF
C11260 sky130_fd_sc_hd__dfrtn_1_8/a_193_47# sky130_fd_sc_hd__dfrtn_1_8/a_448_47# -0.00fF
C11261 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__inv_1_45/Y 0.06fF
C11262 DOUT[13] sky130_fd_sc_hd__dfrtn_1_35/a_1283_21# 0.00fF
C11263 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.00fF
C11264 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__dfrtn_1_26/a_761_289# 0.00fF
C11265 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# 0.00fF
C11266 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# 0.00fF
C11267 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# sky130_fd_sc_hd__dfrtn_1_7/a_27_47# 0.00fF
C11268 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# sky130_fd_sc_hd__dfrtn_1_7/a_193_47# 0.00fF
C11269 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__dfrtn_1_7/a_651_413# 0.00fF
C11270 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__dfrtn_1_7/a_543_47# 0.00fF
C11271 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C11272 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C11273 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_3/a_805_47# 0.00fF
C11274 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_0/a_1217_47# 0.00fF
C11275 sky130_fd_sc_hd__dfrtp_1_0/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11276 sky130_fd_sc_hd__dfrtp_1_0/a_805_47# VDD 0.00fF
C11277 sky130_fd_sc_hd__nand3b_1_0/a_232_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C11278 sky130_fd_sc_hd__nor3_2_3/C out 0.01fF
C11279 sky130_fd_sc_hd__dfrtn_1_21/a_1217_47# RESET_COUNTERn 0.00fF
C11280 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11281 sky130_fd_sc_hd__nor3_1_1/a_109_297# DOUT[5] 0.00fF
C11282 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_48/A 0.01fF
C11283 sky130_fd_sc_hd__nand3b_1_0/a_316_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C11284 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# RESET_COUNTERn 0.12fF
C11285 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# DOUT[7] 0.00fF
C11286 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# DOUT[6] 0.01fF
C11287 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# DOUT[20] 0.00fF
C11288 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C11289 sky130_fd_sc_hd__dfrtn_1_22/a_639_47# RESET_COUNTERn 0.00fF
C11290 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C11291 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C11292 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_805_47# 0.00fF
C11293 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# 0.00fF
C11294 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# 0.00fF
C11295 sky130_fd_sc_hd__dfrtn_1_39/a_1217_47# VDD 0.00fF
C11296 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# 0.01fF
C11297 sky130_fd_sc_hd__dfrtn_1_31/a_543_47# sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C11298 CLK_REF sky130_fd_sc_hd__dfrtn_1_20/a_448_47# 0.00fF
C11299 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C11300 sky130_fd_sc_hd__nor3_1_15/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11301 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# VDD 0.19fF
C11302 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# 0.00fF
C11303 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_10/a_651_413# -0.00fF
C11304 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_10/a_448_47# -0.00fF
C11305 sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# 0.00fF
C11306 sky130_fd_sc_hd__inv_1_32/A DOUT[2] 0.00fF
C11307 sky130_fd_sc_hd__dfrtn_1_14/a_448_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C11308 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# outb 0.00fF
C11309 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C11310 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11311 sky130_fd_sc_hd__dfrtn_1_18/a_1217_47# VDD 0.00fF
C11312 sky130_fd_sc_hd__inv_1_5/A sky130_fd_sc_hd__inv_1_8/Y 0.09fF
C11313 sky130_fd_sc_hd__inv_1_13/A sky130_fd_sc_hd__inv_1_8/A 0.01fF
C11314 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C11315 sky130_fd_sc_hd__dfrtn_1_5/a_805_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C11316 sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# sky130_fd_sc_hd__dfrtn_1_19/a_543_47# 0.00fF
C11317 sky130_fd_sc_hd__dfrtn_1_17/a_1270_413# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C11318 sky130_fd_sc_hd__dfrtn_1_26/a_543_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C11319 sky130_fd_sc_hd__dfrtn_1_16/a_651_413# RESET_COUNTERn 0.00fF
C11320 sky130_fd_sc_hd__dfrtn_1_8/a_1270_413# DOUT[21] 0.00fF
C11321 sky130_fd_sc_hd__dfrtn_1_8/a_543_47# RESET_COUNTERn 0.01fF
C11322 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# DOUT[14] 0.00fF
C11323 sky130_fd_sc_hd__nor3_2_1/a_281_297# out 0.00fF
C11324 VDD sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# 0.00fF
C11325 sky130_fd_sc_hd__dfrtn_1_9/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11326 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# SEL_CONV_TIME[1] 0.01fF
C11327 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__inv_1_30/Y 0.07fF
C11328 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_20/a_651_413# -0.00fF
C11329 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C11330 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# 0.00fF
C11331 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# 0.00fF
C11332 sky130_fd_sc_hd__dfrtn_1_32/a_761_289# sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C11333 sky130_fd_sc_hd__nor3_1_0/a_109_297# DOUT[18] 0.00fF
C11334 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_13/a_193_47# 0.00fF
C11335 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__o2111a_2_0/a_80_21# 0.00fF
C11336 sky130_fd_sc_hd__dfrtn_1_19/a_651_413# VDD 0.01fF
C11337 sky130_fd_sc_hd__dfrtp_1_3/a_805_47# DOUT[23] 0.00fF
C11338 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C11339 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__conb_1_0/LO 0.00fF
C11340 sky130_fd_sc_hd__nor3_1_13/a_193_297# sky130_fd_sc_hd__nor3_1_5/A 0.00fF
C11341 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_1/a_651_413# 0.00fF
C11342 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_1/a_448_47# 0.00fF
C11343 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# sky130_fd_sc_hd__nor3_1_19/Y 0.01fF
C11344 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_18/a_651_413# 0.00fF
C11345 sky130_fd_sc_hd__inv_1_44/Y sky130_fd_sc_hd__o2111a_2_0/X 0.01fF
C11346 sky130_fd_sc_hd__inv_1_41/Y sky130_fd_sc_hd__or3_1_0/C 0.00fF
C11347 sky130_fd_sc_hd__mux4_2_0/a_1281_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C11348 sky130_fd_sc_hd__dfrtn_1_24/a_1462_47# SEL_CONV_TIME[1] 0.00fF
C11349 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# 0.00fF
C11350 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__inv_1_44/Y 0.02fF
C11351 DOUT[4] sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.00fF
C11352 sky130_fd_sc_hd__nor3_1_2/a_109_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11353 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C11354 sky130_fd_sc_hd__or2b_1_0/X sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C11355 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C11356 DOUT[4] sky130_fd_sc_hd__inv_1_9/A 0.01fF
C11357 sky130_fd_sc_hd__dfrtn_1_23/a_805_47# RESET_COUNTERn 0.00fF
C11358 sky130_fd_sc_hd__dfrtn_1_22/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11359 sky130_fd_sc_hd__dfrtn_1_7/a_639_47# DOUT[6] 0.00fF
C11360 sky130_fd_sc_hd__dfrtn_1_7/a_448_47# RESET_COUNTERn 0.00fF
C11361 sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# DOUT[7] 0.00fF
C11362 sky130_fd_sc_hd__dfrtn_1_7/a_805_47# DOUT[20] 0.00fF
C11363 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# 0.00fF
C11364 sky130_fd_sc_hd__dfrtn_1_10/a_805_47# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C11365 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C11366 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# DOUT[3] 0.01fF
C11367 DOUT[4] sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.00fF
C11368 sky130_fd_sc_hd__dfrtn_1_30/a_543_47# sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.00fF
C11369 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_0/a_639_47# -0.00fF
C11370 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C11371 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__dfrtn_1_35/a_193_47# -0.00fF
C11372 sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__inv_1_22/Y 0.00fF
C11373 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# RESET_COUNTERn 0.00fF
C11374 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# CLK_REF 0.01fF
C11375 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__nor2_1_0/a_109_297# 0.00fF
C11376 DOUT[8] RESET_COUNTERn 0.00fF
C11377 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C11378 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C11379 sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C11380 sky130_fd_sc_hd__dfrtn_1_14/a_543_47# DOUT[17] 0.00fF
C11381 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_1290_413# -0.00fF
C11382 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_1478_413# -0.00fF
C11383 sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__mux4_1_0/a_750_97# -0.00fF
C11384 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# sky130_fd_sc_hd__dfrtn_1_27/a_448_47# 0.00fF
C11385 sky130_fd_sc_hd__dfrtn_1_27/a_1270_413# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C11386 sky130_fd_sc_hd__dfrtn_1_26/a_805_47# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C11387 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11388 sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# VDD 0.00fF
C11389 sky130_fd_sc_hd__dfrtn_1_40/a_1270_413# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C11390 sky130_fd_sc_hd__dfrtn_1_16/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C11391 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C11392 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# VDD 0.01fF
C11393 sky130_fd_sc_hd__dfrtn_1_8/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C11394 DOUT[16] sky130_fd_sc_hd__inv_1_36/A 0.00fF
C11395 sky130_fd_sc_hd__dfrtn_1_36/a_193_47# sky130_fd_sc_hd__inv_1_36/A 0.01fF
C11396 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C11397 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_31/a_448_47# 0.00fF
C11398 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C11399 sky130_fd_sc_hd__dfrtn_1_9/a_805_47# DOUT[14] 0.00fF
C11400 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_12/a_761_289# 0.01fF
C11401 DOUT[4] sky130_fd_sc_hd__dfrtn_1_32/a_27_47# 0.01fF
C11402 VDD sky130_fd_sc_hd__inv_1_31/Y 0.13fF
C11403 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_543_47# 0.00fF
C11404 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_761_289# 0.00fF
C11405 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C11406 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C11407 sky130_fd_sc_hd__o211a_1_1/a_510_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C11408 CLK_REF sky130_fd_sc_hd__or2_2_0/a_121_297# 0.00fF
C11409 sky130_fd_sc_hd__or2b_1_0/X sky130_fd_sc_hd__inv_1_49/A 0.03fF
C11410 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_14/a_543_47# 0.00fF
C11411 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__dfrtn_1_14/a_27_47# 0.00fF
C11412 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_14/a_761_289# 0.00fF
C11413 sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# SEL_CONV_TIME[1] 0.00fF
C11414 sky130_fd_sc_hd__dfrtn_1_20/a_1462_47# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C11415 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__dfrtn_1_42/a_27_47# 0.00fF
C11416 sky130_fd_sc_hd__inv_1_4/A DOUT[3] 0.08fF
C11417 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__inv_1_6/A 0.01fF
C11418 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__inv_1_52/A 0.13fF
C11419 sky130_fd_sc_hd__dfrtn_1_23/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11420 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_30/a_1270_413# 0.00fF
C11421 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C11422 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11423 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# VDD 0.05fF
C11424 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# sky130_fd_sc_hd__o221ai_1_0/a_295_297# 0.00fF
C11425 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C11426 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C11427 sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11428 sky130_fd_sc_hd__dfrtn_1_11/a_639_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C11429 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C11430 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_2/A 0.10fF
C11431 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__nor3_1_3/a_109_297# 0.00fF
C11432 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11433 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# VDD 0.00fF
C11434 sky130_fd_sc_hd__inv_1_46/Y SEL_CONV_TIME[1] 0.01fF
C11435 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C11436 sky130_fd_sc_hd__inv_1_18/Y DOUT[10] 0.00fF
C11437 sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# sky130_fd_sc_hd__dfrtn_1_23/a_27_47# 0.00fF
C11438 sky130_fd_sc_hd__dfrtn_1_12/a_761_289# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C11439 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C11440 sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# SEL_CONV_TIME[1] 0.00fF
C11441 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# RESET_COUNTERn 0.01fF
C11442 sky130_fd_sc_hd__inv_1_43/Y RESET_COUNTERn 0.09fF
C11443 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11444 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C11445 sky130_fd_sc_hd__nor2_1_0/a_109_297# DOUT[4] 0.00fF
C11446 sky130_fd_sc_hd__nor3_1_0/a_193_297# RESET_COUNTERn 0.00fF
C11447 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__dfrtn_1_30/a_543_47# 0.00fF
C11448 sky130_fd_sc_hd__nor3_2_3/B DOUT[6] 0.06fF
C11449 sky130_fd_sc_hd__nor3_1_10/a_109_297# DOUT[7] 0.00fF
C11450 sky130_fd_sc_hd__nor3_1_10/a_193_297# DOUT[6] 0.00fF
C11451 sky130_fd_sc_hd__dfrtn_1_33/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C11452 sky130_fd_sc_hd__dfrtn_1_33/a_1108_47# VDD 0.06fF
C11453 sky130_fd_sc_hd__inv_1_9/A outb 0.00fF
C11454 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# RESET_COUNTERn 0.35fF
C11455 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# sky130_fd_sc_hd__inv_1_27/Y 0.00fF
C11456 sky130_fd_sc_hd__dfrtn_1_30/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11457 sky130_fd_sc_hd__dfrtn_1_30/a_805_47# VDD 0.00fF
C11458 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# DOUT[3] 0.00fF
C11459 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C11460 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__nor3_1_4/a_193_297# 0.00fF
C11461 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__nor3_1_4/a_109_297# 0.00fF
C11462 sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# sky130_fd_sc_hd__inv_1_35/A 0.02fF
C11463 sky130_fd_sc_hd__nor3_1_0/a_109_297# DOUT[22] 0.00fF
C11464 DOUT[4] sky130_fd_sc_hd__dfrtn_1_31/a_448_47# 0.00fF
C11465 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C11466 sky130_fd_sc_hd__dfrtn_1_30/a_639_47# sky130_fd_sc_hd__dfrtn_1_31/a_27_47# 0.00fF
C11467 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_639_47# 0.00fF
C11468 sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# sky130_fd_sc_hd__dfrtn_1_28/a_27_47# 0.00fF
C11469 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C11470 sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# DOUT[14] 0.00fF
C11471 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C11472 sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C11473 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C11474 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__dfrtn_1_17/a_651_413# 0.00fF
C11475 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# HEADER_0/a_508_138# 0.00fF
C11476 sky130_fd_sc_hd__inv_1_42/A DOUT[21] 0.12fF
C11477 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# DOUT[17] 0.01fF
C11478 sky130_fd_sc_hd__dfrtn_1_34/a_651_413# SEL_CONV_TIME[1] 0.00fF
C11479 sky130_fd_sc_hd__o211a_1_1/a_297_297# sky130_fd_sc_hd__dfrtn_1_17/a_651_413# 0.00fF
C11480 sky130_fd_sc_hd__nor3_1_14/a_109_297# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C11481 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C11482 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# sky130_fd_sc_hd__dfrtn_1_29/a_761_289# 0.00fF
C11483 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# sky130_fd_sc_hd__dfrtn_1_29/a_543_47# 0.00fF
C11484 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# 0.00fF
C11485 sky130_fd_sc_hd__dfrtn_1_25/a_639_47# SEL_CONV_TIME[0] 0.00fF
C11486 sky130_fd_sc_hd__nand3b_1_1/a_316_47# DOUT[21] 0.00fF
C11487 sky130_fd_sc_hd__or3_1_0/a_183_297# DOUT[21] 0.00fF
C11488 sky130_fd_sc_hd__dfrtn_1_38/a_543_47# VDD 0.04fF
C11489 sky130_fd_sc_hd__dfrtn_1_36/a_1462_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C11490 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# 0.00fF
C11491 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# 0.00fF
C11492 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# sky130_fd_sc_hd__inv_1_45/A 0.31fF
C11493 sky130_fd_sc_hd__nor3_1_6/a_193_297# DOUT[9] 0.00fF
C11494 sky130_fd_sc_hd__or3b_2_0/B DONE 0.01fF
C11495 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_11/a_1270_413# 0.00fF
C11496 sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# 0.00fF
C11497 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# sky130_fd_sc_hd__dfrtn_1_11/a_761_289# 0.00fF
C11498 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__dfrtn_1_11/a_543_47# 0.00fF
C11499 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_639_47# 0.00fF
C11500 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C11501 sky130_fd_sc_hd__dfrtn_1_42/a_193_47# DOUT[15] 0.00fF
C11502 DOUT[4] sky130_fd_sc_hd__dfrtn_1_32/a_1217_47# 0.00fF
C11503 DOUT[12] sky130_fd_sc_hd__inv_1_8/A 0.01fF
C11504 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# -0.00fF
C11505 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_1/a_448_47# -0.00fF
C11506 sky130_fd_sc_hd__dfrtn_1_12/a_805_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C11507 sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# sky130_fd_sc_hd__inv_1_6/A 0.02fF
C11508 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__dfrtn_1_40/a_1270_413# 0.00fF
C11509 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__dfrtn_1_17/a_651_413# 0.00fF
C11510 sky130_fd_sc_hd__dfrtn_1_12/a_805_47# sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# 0.00fF
C11511 sky130_fd_sc_hd__dfrtn_1_12/a_639_47# sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# 0.00fF
C11512 sky130_fd_sc_hd__dfrtn_1_12/a_761_289# sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# 0.00fF
C11513 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# 0.00fF
C11514 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# sky130_fd_sc_hd__dfrtn_1_37/a_543_47# -0.00fF
C11515 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# -0.00fF
C11516 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# -0.00fF
C11517 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# 0.00fF
C11518 sky130_fd_sc_hd__dfrtn_1_28/a_448_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C11519 sky130_fd_sc_hd__dfrtn_1_26/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11520 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11521 sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# VDD 0.05fF
C11522 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C11523 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# DOUT[14] 0.00fF
C11524 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C11525 sky130_fd_sc_hd__or3_1_0/a_183_297# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C11526 sky130_fd_sc_hd__inv_1_6/A DOUT[7] 0.08fF
C11527 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C11528 sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11529 sky130_fd_sc_hd__dfrtn_1_34/a_448_47# VDD 0.01fF
C11530 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_7/a_543_47# 0.00fF
C11531 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# 0.00fF
C11532 sky130_fd_sc_hd__or2b_1_0/a_301_297# sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# 0.00fF
C11533 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_8/a_27_47# 0.01fF
C11534 sky130_fd_sc_hd__dfrtn_1_29/a_805_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C11535 sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C11536 sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# sky130_fd_sc_hd__inv_1_40/Y 0.01fF
C11537 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_543_47# -0.00fF
C11538 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_3/a_761_289# -0.00fF
C11539 sky130_fd_sc_hd__dfrtn_1_28/a_448_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C11540 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C11541 sky130_fd_sc_hd__o2111a_2_0/a_458_47# SEL_CONV_TIME[1] 0.00fF
C11542 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# RESET_COUNTERn 0.01fF
C11543 sky130_fd_sc_hd__dfrtn_1_25/a_1270_413# DOUT[21] 0.00fF
C11544 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11545 DOUT[23] lc_out 0.00fF
C11546 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_6/a_639_47# 0.00fF
C11547 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__nor3_2_3/B 0.11fF
C11548 sky130_fd_sc_hd__dfrtp_1_1/a_805_47# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C11549 sky130_fd_sc_hd__inv_1_4/A DOUT[20] 0.01fF
C11550 sky130_fd_sc_hd__dfrtn_1_25/a_1462_47# sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C11551 sky130_fd_sc_hd__dfrtn_1_32/a_1270_413# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C11552 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C11553 sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C11554 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C11555 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.01fF
C11556 DOUT[9] sky130_fd_sc_hd__dfrtn_1_6/a_448_47# 0.00fF
C11557 sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# DOUT[3] 0.00fF
C11558 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# DOUT[15] 0.00fF
C11559 sky130_fd_sc_hd__dfrtn_1_3/a_1462_47# RESET_COUNTERn 0.00fF
C11560 sky130_fd_sc_hd__or3b_2_0/a_472_297# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C11561 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.01fF
C11562 sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C11563 DOUT[19] DOUT[14] 0.04fF
C11564 DOUT[4] sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C11565 DOUT[13] sky130_fd_sc_hd__or3b_2_0/a_27_47# 0.00fF
C11566 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__inv_1_43/A 0.01fF
C11567 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# 0.00fF
C11568 sky130_fd_sc_hd__dfrtn_1_7/a_448_47# HEADER_0/a_508_138# 0.00fF
C11569 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11570 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# SEL_CONV_TIME[1] 0.00fF
C11571 sky130_fd_sc_hd__nor3_1_4/A sky130_fd_sc_hd__inv_1_13/A 0.00fF
C11572 sky130_fd_sc_hd__inv_1_13/Y sky130_fd_sc_hd__inv_1_5/Y 0.02fF
C11573 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# VDD 0.00fF
C11574 sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# RESET_COUNTERn 0.03fF
C11575 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__inv_1_44/A 0.02fF
C11576 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# SEL_CONV_TIME[3] 0.00fF
C11577 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C11578 sky130_fd_sc_hd__nor3_1_12/a_109_297# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C11579 sky130_fd_sc_hd__dfrtn_1_0/a_1217_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C11580 sky130_fd_sc_hd__nor3_1_16/a_109_297# RESET_COUNTERn 0.00fF
C11581 sky130_fd_sc_hd__dfrtn_1_11/a_761_289# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C11582 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_10/a_1283_21# 0.00fF
C11583 sky130_fd_sc_hd__dfrtn_1_0/a_1270_413# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C11584 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C11585 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C11586 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtp_1_3/a_761_289# 0.00fF
C11587 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtp_1_3/a_448_47# 0.00fF
C11588 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__mux4_2_0/a_288_47# -0.00fF
C11589 sky130_fd_sc_hd__dfrtp_1_1/a_805_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C11590 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C11591 HEADER_0/a_508_138# DOUT[8] 0.00fF
C11592 sky130_fd_sc_hd__dfrtn_1_0/a_1217_47# DOUT[17] 0.00fF
C11593 sky130_fd_sc_hd__o2111a_2_0/a_386_47# VDD 0.00fF
C11594 sky130_fd_sc_hd__inv_1_24/A DOUT[12] 0.00fF
C11595 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# sky130_fd_sc_hd__dfrtn_1_29/a_651_413# 0.00fF
C11596 sky130_fd_sc_hd__dfrtn_1_24/a_651_413# sky130_fd_sc_hd__dfrtn_1_29/a_639_47# 0.00fF
C11597 sky130_fd_sc_hd__dfrtn_1_17/a_1270_413# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C11598 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# DOUT[20] 0.00fF
C11599 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# DOUT[8] 0.00fF
C11600 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# RESET_COUNTERn 0.02fF
C11601 sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C11602 sky130_fd_sc_hd__dfrtn_1_4/a_1270_413# RESET_COUNTERn -0.00fF
C11603 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# SEL_CONV_TIME[0] 0.00fF
C11604 sky130_fd_sc_hd__dfrtn_1_38/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11605 sky130_fd_sc_hd__dfrtn_1_33/a_1462_47# sky130_fd_sc_hd__inv_1_45/A 0.00fF
C11606 DOUT[13] sky130_fd_sc_hd__nor3_2_3/C 0.06fF
C11607 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__dfrtn_1_34/a_193_47# 0.00fF
C11608 sky130_fd_sc_hd__or2b_1_0/a_301_297# sky130_fd_sc_hd__dfrtn_1_34/a_27_47# 0.00fF
C11609 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__nor3_1_3/a_193_297# 0.00fF
C11610 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__nor3_1_3/a_109_297# 0.00fF
C11611 sky130_fd_sc_hd__nor3_1_19/a_193_297# VDD 0.00fF
C11612 SLC_0/a_438_293# RESET_COUNTERn 0.01fF
C11613 sky130_fd_sc_hd__dfrtn_1_42/a_1462_47# DOUT[15] 0.00fF
C11614 sky130_fd_sc_hd__dfrtn_1_31/a_543_47# sky130_fd_sc_hd__inv_1_49/A 0.02fF
C11615 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# 0.00fF
C11616 DOUT[13] sky130_fd_sc_hd__dfrtn_1_31/a_193_47# 0.02fF
C11617 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# SEL_CONV_TIME[2] 0.01fF
C11618 SEL_CONV_TIME[1] sky130_fd_sc_hd__mux4_1_0/X 0.02fF
C11619 DOUT[23] sky130_fd_sc_hd__nor3_2_3/B 0.04fF
C11620 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_8/A 0.31fF
C11621 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.26fF
C11622 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__o2111a_2_0/X 0.01fF
C11623 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C11624 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.04fF
C11625 sky130_fd_sc_hd__dfrtn_1_14/a_448_47# VDD 0.00fF
C11626 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__dfrtn_1_0/a_651_413# 0.00fF
C11627 sky130_fd_sc_hd__dfrtn_1_12/a_651_413# sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# 0.00fF
C11628 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C11629 sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11630 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# 0.00fF
C11631 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C11632 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# RESET_COUNTERn 0.00fF
C11633 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__inv_1_22/A 0.34fF
C11634 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__inv_1_8/Y 0.01fF
C11635 VDD sky130_fd_sc_hd__inv_1_5/A 0.28fF
C11636 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__inv_1_45/Y 0.01fF
C11637 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C11638 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_41/a_805_47# -0.00fF
C11639 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__dfrtn_1_41/a_639_47# -0.00fF
C11640 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C11641 sky130_fd_sc_hd__inv_1_50/Y RESET_COUNTERn 0.01fF
C11642 sky130_fd_sc_hd__dfrtn_1_3/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11643 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_8/a_1217_47# 0.00fF
C11644 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# sky130_fd_sc_hd__inv_1_2/A 0.01fF
C11645 sky130_fd_sc_hd__dfrtn_1_39/a_651_413# RESET_COUNTERn 0.00fF
C11646 sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C11647 sky130_fd_sc_hd__dfrtn_1_22/a_1108_47# sky130_fd_sc_hd__inv_1_39/Y 0.03fF
C11648 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C11649 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__inv_1_13/A 0.02fF
C11650 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# DOUT[21] 0.02fF
C11651 sky130_fd_sc_hd__dfrtn_1_42/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C11652 sky130_fd_sc_hd__dfrtp_1_3/a_805_47# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C11653 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__inv_1_48/A 0.00fF
C11654 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__nor3_1_3/a_109_297# 0.00fF
C11655 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__nor3_1_3/a_193_297# 0.00fF
C11656 sky130_fd_sc_hd__dfrtn_1_37/a_805_47# sky130_fd_sc_hd__inv_1_32/Y 0.00fF
C11657 DOUT[9] sky130_fd_sc_hd__nor3_1_1/a_193_297# 0.00fF
C11658 sky130_fd_sc_hd__dfrtn_1_18/a_651_413# RESET_COUNTERn -0.00fF
C11659 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__dfrtn_1_25/a_193_47# 0.00fF
C11660 sky130_fd_sc_hd__or3_1_0/a_111_297# sky130_fd_sc_hd__dfrtn_1_25/a_27_47# 0.00fF
C11661 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# 0.00fF
C11662 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# 0.00fF
C11663 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C11664 DOUT[4] sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# 0.00fF
C11665 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C11666 sky130_fd_sc_hd__dfrtn_1_4/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11667 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# SEL_CONV_TIME[0] 0.03fF
C11668 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# SEL_CONV_TIME[3] 0.00fF
C11669 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C11670 sky130_fd_sc_hd__inv_1_14/A DOUT[22] 0.00fF
C11671 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__dfrtn_1_7/a_27_47# 0.00fF
C11672 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# DOUT[3] 0.01fF
C11673 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# VDD 0.05fF
C11674 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C11675 sky130_fd_sc_hd__mux4_2_0/a_1279_413# sky130_fd_sc_hd__o311a_1_0/a_266_47# 0.00fF
C11676 sky130_fd_sc_hd__mux4_2_0/a_1281_47# sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.00fF
C11677 sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# RESET_COUNTERn 0.04fF
C11678 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_27_47# 0.00fF
C11679 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__mux4_2_0/a_1279_413# -0.00fF
C11680 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C11681 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# 0.00fF
C11682 sky130_fd_sc_hd__dfrtn_1_19/a_543_47# RESET_COUNTERn 0.02fF
C11683 sky130_fd_sc_hd__dfrtn_1_41/a_651_413# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C11684 CLK_REF sky130_fd_sc_hd__dfrtn_1_17/a_651_413# 0.00fF
C11685 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C11686 sky130_fd_sc_hd__o311a_1_0/a_81_21# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C11687 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C11688 sky130_fd_sc_hd__dfrtp_1_0/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11689 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C11690 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_543_47# 0.00fF
C11691 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_761_289# 0.00fF
C11692 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C11693 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C11694 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__inv_1_8/A 0.02fF
C11695 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_448_47# -0.00fF
C11696 sky130_fd_sc_hd__dfrtn_1_21/a_1217_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C11697 sky130_fd_sc_hd__or3b_2_0/a_388_297# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C11698 sky130_fd_sc_hd__dfrtn_1_35/a_543_47# sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.00fF
C11699 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_651_413# 0.00fF
C11700 sky130_fd_sc_hd__dfrtn_1_35/a_761_289# sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# 0.00fF
C11701 sky130_fd_sc_hd__dfrtn_1_35/a_448_47# sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C11702 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_25/a_651_413# -0.00fF
C11703 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__dfrtn_1_25/a_448_47# -0.00fF
C11704 DOUT[13] sky130_fd_sc_hd__dfrtn_1_31/a_1462_47# 0.00fF
C11705 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# 0.00fF
C11706 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_805_47# 0.00fF
C11707 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__inv_1_7/Y 0.01fF
C11708 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C11709 sky130_fd_sc_hd__dfrtn_1_28/a_805_47# VDD 0.00fF
C11710 sky130_fd_sc_hd__dfrtn_1_23/a_448_47# sky130_fd_sc_hd__inv_1_39/Y 0.00fF
C11711 sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C11712 DOUT[4] sky130_fd_sc_hd__inv_1_51/Y 0.03fF
C11713 DOUT[1] sky130_fd_sc_hd__inv_1_40/A 0.48fF
C11714 sky130_fd_sc_hd__dfrtn_1_4/a_1270_413# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C11715 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# sky130_fd_sc_hd__inv_1_43/A 0.03fF
C11716 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__inv_1_5/A 0.01fF
C11717 sky130_fd_sc_hd__dfrtn_1_25/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11718 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# 0.02fF
C11719 sky130_fd_sc_hd__dfrtn_1_12/a_761_289# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C11720 sky130_fd_sc_hd__dfrtn_1_9/a_448_47# sky130_fd_sc_hd__inv_1_12/A 0.02fF
C11721 sky130_fd_sc_hd__dfrtn_1_0/a_543_47# VDD 0.06fF
C11722 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11723 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11724 sky130_fd_sc_hd__dfrtn_1_16/a_651_413# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C11725 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C11726 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__inv_1_14/A 0.01fF
C11727 sky130_fd_sc_hd__mux4_1_0/a_193_47# SEL_CONV_TIME[1] 0.00fF
C11728 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C11729 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_38/a_651_413# 0.00fF
C11730 DOUT[9] sky130_fd_sc_hd__dfrtn_1_3/a_448_47# 0.00fF
C11731 sky130_fd_sc_hd__nor3_1_3/a_109_297# VIN 0.00fF
C11732 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C11733 VDD sky130_fd_sc_hd__nor3_1_5/a_193_297# 0.00fF
C11734 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_14/a_761_289# 0.01fF
C11735 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C11736 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C11737 sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# sky130_fd_sc_hd__inv_1_32/Y 0.00fF
C11738 sky130_fd_sc_hd__dfrtn_1_20/a_1270_413# VDD 0.00fF
C11739 sky130_fd_sc_hd__dfrtn_1_24/a_1462_47# DOUT[21] 0.00fF
C11740 sky130_fd_sc_hd__dfrtn_1_24/a_651_413# RESET_COUNTERn 0.00fF
C11741 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# DOUT[20] 0.00fF
C11742 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# RESET_COUNTERn 0.03fF
C11743 sky130_fd_sc_hd__dfrtn_1_25/a_805_47# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C11744 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C11745 sky130_fd_sc_hd__dfrtn_1_9/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11746 sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# sky130_fd_sc_hd__inv_1_32/Y 0.01fF
C11747 sky130_fd_sc_hd__dfrtp_1_3/a_1217_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C11748 DOUT[1] sky130_fd_sc_hd__dfrtn_1_36/a_1270_413# 0.00fF
C11749 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_2/a_761_289# 0.01fF
C11750 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# outb 0.00fF
C11751 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C11752 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__inv_1_31/A 0.00fF
C11753 sky130_fd_sc_hd__dfrtn_1_23/a_805_47# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C11754 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_26/a_639_47# 0.00fF
C11755 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_12/a_761_289# -0.00fF
C11756 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C11757 sky130_fd_sc_hd__dfrtn_1_16/a_1108_47# DOUT[2] 0.01fF
C11758 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# sky130_fd_sc_hd__dfrtn_1_42/a_639_47# -0.00fF
C11759 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__dfrtn_1_13/a_27_47# 0.00fF
C11760 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_761_289# 0.00fF
C11761 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_543_47# 0.00fF
C11762 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# sky130_fd_sc_hd__dfrtn_1_13/a_193_47# 0.00fF
C11763 sky130_fd_sc_hd__o221ai_1_0/a_109_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11764 DOUT[9] sky130_fd_sc_hd__dfrtn_1_4/a_761_289# 0.00fF
C11765 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# DOUT[11] 0.00fF
C11766 sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# SEL_CONV_TIME[0] 0.00fF
C11767 DOUT[1] VDD 4.69fF
C11768 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C11769 sky130_fd_sc_hd__mux4_1_0/a_27_47# VDD 0.01fF
C11770 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C11771 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__inv_1_4/Y 0.01fF
C11772 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C11773 sky130_fd_sc_hd__nor3_2_1/A VDD 0.29fF
C11774 sky130_fd_sc_hd__dfrtn_1_10/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11775 sky130_fd_sc_hd__o211a_1_0/a_79_21# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C11776 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_19/a_448_47# 0.00fF
C11777 sky130_fd_sc_hd__o211a_1_0/a_215_47# VDD 0.00fF
C11778 sky130_fd_sc_hd__inv_1_33/A sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11779 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# VIN 0.04fF
C11780 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# 0.00fF
C11781 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C11782 sky130_fd_sc_hd__dfrtp_1_0/a_639_47# DOUT[23] 0.00fF
C11783 sky130_fd_sc_hd__dfrtn_1_24/a_1462_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C11784 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# 0.01fF
C11785 DOUT[23] DOUT[0] 0.03fF
C11786 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_651_413# -0.00fF
C11787 sky130_fd_sc_hd__dfrtn_1_27/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_448_47# -0.00fF
C11788 sky130_fd_sc_hd__nor3_1_13/a_109_297# DOUT[21] 0.00fF
C11789 sky130_fd_sc_hd__nor3_1_15/a_193_297# DOUT[13] 0.00fF
C11790 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C11791 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_11/a_448_47# 0.00fF
C11792 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C11793 sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# SEL_CONV_TIME[0] 0.00fF
C11794 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# -0.00fF
C11795 sky130_fd_sc_hd__mux4_2_0/a_397_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C11796 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# DOUT[7] 0.00fF
C11797 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# DOUT[6] 0.00fF
C11798 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# RESET_COUNTERn 0.02fF
C11799 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_4/a_639_47# 0.00fF
C11800 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_4/a_805_47# 0.00fF
C11801 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__dfrtn_1_4/a_651_413# 0.00fF
C11802 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__dfrtn_1_4/a_448_47# 0.00fF
C11803 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__dfrtn_1_4/a_543_47# 0.00fF
C11804 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# sky130_fd_sc_hd__dfrtn_1_4/a_761_289# 0.00fF
C11805 sky130_fd_sc_hd__dfrtn_1_39/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_543_47# -0.00fF
C11806 sky130_fd_sc_hd__dfrtn_1_39/a_651_413# SEL_CONV_TIME[2] 0.00fF
C11807 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_38/A 0.00fF
C11808 VDD sky130_fd_sc_hd__or2_2_0/B 0.85fF
C11809 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__o311a_1_0/a_266_47# 0.00fF
C11810 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__o311a_1_0/a_585_47# 0.00fF
C11811 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__o311a_1_0/a_368_297# 0.00fF
C11812 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__inv_1_45/A 0.00fF
C11813 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.01fF
C11814 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# RESET_COUNTERn -0.01fF
C11815 DOUT[1] sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# 0.00fF
C11816 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# DOUT[19] 0.00fF
C11817 sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C11818 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C11819 sky130_fd_sc_hd__dfrtn_1_27/a_1217_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C11820 sky130_fd_sc_hd__nor3_1_1/a_109_297# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C11821 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C11822 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__mux4_2_0/a_600_345# 0.00fF
C11823 sky130_fd_sc_hd__dfrtn_1_35/a_805_47# VDD 0.00fF
C11824 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C11825 sky130_fd_sc_hd__dfrtn_1_30/a_448_47# RESET_COUNTERn 0.00fF
C11826 sky130_fd_sc_hd__dfrtn_1_12/a_805_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C11827 sky130_fd_sc_hd__dfrtn_1_21/a_193_47# sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# -0.00fF
C11828 SLC_0/a_438_293# SLC_0/a_264_22# -0.00fF
C11829 sky130_fd_sc_hd__nor3_2_1/a_27_297# sky130_fd_sc_hd__o211a_1_0/a_297_297# 0.00fF
C11830 sky130_fd_sc_hd__nor3_2_1/a_281_297# sky130_fd_sc_hd__o211a_1_0/a_79_21# 0.00fF
C11831 SLC_0/a_919_243# sky130_fd_sc_hd__inv_1_26/A 0.01fF
C11832 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C11833 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.00fF
C11834 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C11835 sky130_fd_sc_hd__dfrtn_1_18/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# -0.00fF
C11836 sky130_fd_sc_hd__dfrtn_1_18/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_543_47# -0.00fF
C11837 sky130_fd_sc_hd__dfrtn_1_26/a_651_413# SEL_CONV_TIME[0] 0.00fF
C11838 sky130_fd_sc_hd__mux4_2_0/a_193_47# SEL_CONV_TIME[1] -0.00fF
C11839 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# DOUT[19] 0.00fF
C11840 sky130_fd_sc_hd__dfrtn_1_27/a_639_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C11841 sky130_fd_sc_hd__dfrtn_1_34/a_1270_413# SEL_CONV_TIME[0] 0.00fF
C11842 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11843 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# VDD 0.01fF
C11844 sky130_fd_sc_hd__dfrtn_1_23/a_1217_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C11845 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_30/a_1270_413# 0.00fF
C11846 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C11847 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C11848 sky130_fd_sc_hd__inv_1_0/A DOUT[18] 0.01fF
C11849 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C11850 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__nor3_1_4/A 0.03fF
C11851 sky130_fd_sc_hd__inv_1_46/Y DOUT[21] 0.00fF
C11852 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C11853 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C11854 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# -0.00fF
C11855 sky130_fd_sc_hd__dfrtp_1_0/a_1283_21# SLC_0/a_1235_416# 0.00fF
C11856 sky130_fd_sc_hd__dfrtp_1_0/a_1108_47# SLC_0/a_919_243# 0.00fF
C11857 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# SLC_0/a_264_22# 0.00fF
C11858 sky130_fd_sc_hd__dfrtn_1_16/a_761_289# sky130_fd_sc_hd__inv_1_25/A 0.00fF
C11859 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# SLC_0/a_438_293# 0.00fF
C11860 sky130_fd_sc_hd__dfrtp_1_0/a_1270_413# sky130_fd_sc_hd__inv_1_26/A 0.00fF
C11861 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# DOUT[18] 0.00fF
C11862 sky130_fd_sc_hd__inv_1_26/A out 0.01fF
C11863 CLK_REF sky130_fd_sc_hd__dfrtp_1_3/a_805_47# 0.00fF
C11864 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__inv_1_7/A 0.00fF
C11865 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# 0.00fF
C11866 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# 0.01fF
C11867 sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C11868 outb DOUT[15] 0.00fF
C11869 sky130_fd_sc_hd__dfrtn_1_8/a_651_413# outb 0.00fF
C11870 sky130_fd_sc_hd__o211a_1_1/a_510_47# RESET_COUNTERn 0.00fF
C11871 sky130_fd_sc_hd__nor3_2_2/a_281_297# sky130_fd_sc_hd__inv_1_25/A 0.02fF
C11872 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_10/a_761_289# 0.03fF
C11873 sky130_fd_sc_hd__inv_1_36/A RESET_COUNTERn 0.24fF
C11874 sky130_fd_sc_hd__dfrtn_1_10/a_639_47# sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# 0.00fF
C11875 sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# VIN 0.00fF
C11876 sky130_fd_sc_hd__o311a_1_0/a_585_47# VDD 0.00fF
C11877 sky130_fd_sc_hd__o311a_1_0/a_368_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11878 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_12/a_651_413# 0.00fF
C11879 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C11880 sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C11881 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C11882 sky130_fd_sc_hd__mux4_2_0/a_372_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11883 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C11884 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.64fF
C11885 sky130_fd_sc_hd__mux4_2_0/a_600_345# VDD 0.04fF
C11886 sky130_fd_sc_hd__dfrtp_1_0/a_1108_47# out 0.00fF
C11887 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_5/A 0.00fF
C11888 sky130_fd_sc_hd__inv_1_4/Y DOUT[8] 0.01fF
C11889 sky130_fd_sc_hd__inv_1_1/A DOUT[18] 0.01fF
C11890 sky130_fd_sc_hd__dfrtn_1_27/a_543_47# SEL_CONV_TIME[1] 0.00fF
C11891 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# RESET_COUNTERn 0.36fF
C11892 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_2/a_193_47# 0.02fF
C11893 sky130_fd_sc_hd__dfrtn_1_34/a_805_47# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C11894 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C11895 sky130_fd_sc_hd__inv_1_53/A sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C11896 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__nor3_1_4/A 0.22fF
C11897 sky130_fd_sc_hd__dfrtp_1_1/a_448_47# sky130_fd_sc_hd__nor3_2_1/a_27_297# 0.00fF
C11898 sky130_fd_sc_hd__dfrtn_1_33/a_761_289# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C11899 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C11900 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__nand2_1_1/a_113_47# 0.00fF
C11901 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.02fF
C11902 sky130_fd_sc_hd__o2111a_2_0/a_566_47# SEL_CONV_TIME[0] 0.00fF
C11903 sky130_fd_sc_hd__dfrtn_1_35/a_1108_47# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C11904 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# sky130_fd_sc_hd__nor3_2_3/A 0.55fF
C11905 sky130_fd_sc_hd__dfrtn_1_11/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11906 sky130_fd_sc_hd__inv_1_41/Y RESET_COUNTERn 0.00fF
C11907 sky130_fd_sc_hd__dfrtn_1_34/a_651_413# DOUT[21] 0.00fF
C11908 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# RESET_COUNTERn 0.00fF
C11909 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__nand2_1_2/Y 0.00fF
C11910 sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# VDD 0.09fF
C11911 sky130_fd_sc_hd__dfrtp_1_2/a_639_47# RESET_COUNTERn 0.00fF
C11912 sky130_fd_sc_hd__dfrtn_1_35/a_1283_21# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C11913 sky130_fd_sc_hd__dfrtn_1_17/a_1462_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C11914 sky130_fd_sc_hd__nor3_1_20/a_109_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11915 HEADER_1/a_508_138# DOUT[11] 0.02fF
C11916 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__inv_1_33/A 0.00fF
C11917 sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11918 sky130_fd_sc_hd__dfrtn_1_41/a_639_47# VDD 0.00fF
C11919 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C11920 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# DOUT[2] 0.00fF
C11921 sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C11922 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# 0.00fF
C11923 sky130_fd_sc_hd__dfrtn_1_8/a_761_289# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C11924 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_39/a_805_47# 0.00fF
C11925 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# DONE 0.00fF
C11926 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.04fF
C11927 sky130_fd_sc_hd__nor3_1_11/a_193_297# DOUT[14] 0.00fF
C11928 DOUT[9] sky130_fd_sc_hd__inv_1_2/Y 0.01fF
C11929 sky130_fd_sc_hd__nor3_1_4/a_193_297# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C11930 sky130_fd_sc_hd__dfrtn_1_33/a_1462_47# RESET_COUNTERn 0.00fF
C11931 sky130_fd_sc_hd__dfrtn_1_7/a_1462_47# DOUT[19] 0.00fF
C11932 sky130_fd_sc_hd__dfrtn_1_28/a_193_47# SEL_CONV_TIME[0] 0.00fF
C11933 sky130_fd_sc_hd__mux4_2_0/a_872_316# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C11934 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_15/A 0.07fF
C11935 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11936 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C11937 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C11938 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C11939 sky130_fd_sc_hd__dfrtn_1_27/a_761_289# VDD 0.05fF
C11940 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# 0.00fF
C11941 sky130_fd_sc_hd__dfrtn_1_34/a_651_413# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C11942 sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__o211a_1_0/X 0.02fF
C11943 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_18/a_761_289# 0.01fF
C11944 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__dfrtn_1_1/a_193_47# 0.00fF
C11945 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__dfrtn_1_1/a_27_47# 0.00fF
C11946 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# RESET_COUNTERn 0.01fF
C11947 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C11948 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__dfrtp_1_1/D 0.00fF
C11949 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__inv_1_45/Y 0.01fF
C11950 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__inv_1_45/A 0.00fF
C11951 sky130_fd_sc_hd__o211a_1_1/a_297_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11952 sky130_fd_sc_hd__dfrtn_1_37/a_805_47# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C11953 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_761_289# -0.00fF
C11954 sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C11955 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11956 sky130_fd_sc_hd__o2111a_2_0/a_458_47# DOUT[21] 0.00fF
C11957 sky130_fd_sc_hd__o221ai_1_0/a_213_123# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C11958 sky130_fd_sc_hd__o2111a_2_0/X sky130_fd_sc_hd__nor3_2_3/B 0.03fF
C11959 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C11960 sky130_fd_sc_hd__or3b_2_0/a_472_297# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C11961 sky130_fd_sc_hd__dfrtn_1_38/a_805_47# RESET_COUNTERn 0.00fF
C11962 sky130_fd_sc_hd__dfrtn_1_26/a_761_289# sky130_fd_sc_hd__inv_1_43/Y 0.01fF
C11963 sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C11964 sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# DOUT[18] 0.00fF
C11965 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_21/a_651_413# 0.00fF
C11966 sky130_fd_sc_hd__inv_1_49/A RESET_COUNTERn 0.98fF
C11967 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11968 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# VDD 0.08fF
C11969 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__inv_1_4/A 0.00fF
C11970 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C11971 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_448_47# 0.00fF
C11972 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C11973 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C11974 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C11975 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.00fF
C11976 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11977 sky130_fd_sc_hd__nor3_1_10/a_109_297# VIN 0.00fF
C11978 sky130_fd_sc_hd__dfrtp_1_3/a_1283_21# sky130_fd_sc_hd__or2_2_0/B 0.02fF
C11979 sky130_fd_sc_hd__inv_1_10/A DOUT[1] 0.01fF
C11980 sky130_fd_sc_hd__or2_2_0/B sky130_fd_sc_hd__o211a_1_0/X 0.00fF
C11981 sky130_fd_sc_hd__nand2_1_2/Y DOUT[4] 0.01fF
C11982 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.64fF
C11983 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# VDD 0.07fF
C11984 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C11985 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__inv_1_44/A 0.01fF
C11986 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_30/a_543_47# 0.00fF
C11987 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11988 sky130_fd_sc_hd__dfrtn_1_39/a_805_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C11989 sky130_fd_sc_hd__dfrtn_1_17/a_448_47# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C11990 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# DOUT[21] 0.02fF
C11991 sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# DOUT[23] 0.00fF
C11992 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C11993 DOUT[13] sky130_fd_sc_hd__inv_1_50/A 0.01fF
C11994 sky130_fd_sc_hd__dfrtn_1_0/a_543_47# DOUT[5] 0.00fF
C11995 sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C11996 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_639_47# -0.00fF
C11997 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# DOUT[14] 0.00fF
C11998 sky130_fd_sc_hd__mux4_1_0/a_27_413# SEL_CONV_TIME[0] 0.00fF
C11999 sky130_fd_sc_hd__dfrtn_1_14/a_761_289# RESET_COUNTERn 0.02fF
C12000 sky130_fd_sc_hd__dfrtn_1_28/a_1283_21# sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C12001 sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# sky130_fd_sc_hd__dfrtn_1_13/a_193_47# 0.00fF
C12002 sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# sky130_fd_sc_hd__dfrtn_1_13/a_27_47# 0.00fF
C12003 sky130_fd_sc_hd__o2111a_2_0/a_458_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C12004 sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# sky130_fd_sc_hd__nor3_2_2/A 0.01fF
C12005 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__inv_1_47/Y 0.00fF
C12006 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# 0.00fF
C12007 sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# RESET_COUNTERn 0.00fF
C12008 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# 0.01fF
C12009 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C12010 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C12011 sky130_fd_sc_hd__inv_1_0/A DOUT[22] 0.00fF
C12012 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_44/Y 0.01fF
C12013 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# sky130_fd_sc_hd__dfrtp_1_3/a_651_413# 0.00fF
C12014 sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# sky130_fd_sc_hd__dfrtp_1_3/a_543_47# 0.00fF
C12015 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__dfrtp_1_3/a_639_47# 0.00fF
C12016 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_805_47# 0.00fF
C12017 sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C12018 sky130_fd_sc_hd__dfrtp_1_1/a_805_47# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C12019 DOUT[23] DOUT[2] 0.02fF
C12020 DOUT[15] sky130_fd_sc_hd__nor3_2_3/A 0.19fF
C12021 sky130_fd_sc_hd__dfrtn_1_16/a_1217_47# sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C12022 sky130_fd_sc_hd__dfrtn_1_20/a_543_47# sky130_fd_sc_hd__dfrtn_1_21/a_761_289# 0.00fF
C12023 sky130_fd_sc_hd__dfrtn_1_33/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12024 sky130_fd_sc_hd__nor3_1_5/a_193_297# DOUT[5] 0.00fF
C12025 sky130_fd_sc_hd__dfrtn_1_19/a_193_47# sky130_fd_sc_hd__dfrtn_1_19/a_448_47# -0.00fF
C12026 sky130_fd_sc_hd__dfrtn_1_19/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_651_413# -0.00fF
C12027 sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# sky130_fd_sc_hd__inv_1_40/A 0.00fF
C12028 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C12029 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__nand3b_1_1/a_53_93# 0.00fF
C12030 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# DOUT[22] 0.00fF
C12031 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__dfrtn_1_34/a_27_47# 0.00fF
C12032 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# 0.01fF
C12033 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_37/a_651_413# 0.00fF
C12034 sky130_fd_sc_hd__dfrtn_1_40/a_1270_413# sky130_fd_sc_hd__dfrtn_1_37/a_27_47# 0.00fF
C12035 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__dfrtn_1_37/a_543_47# 0.00fF
C12036 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_37/a_193_47# 0.00fF
C12037 sky130_fd_sc_hd__dfrtn_1_24/a_448_47# sky130_fd_sc_hd__inv_1_48/A 0.01fF
C12038 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C12039 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C12040 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C12041 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_651_413# 0.00fF
C12042 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# 0.00fF
C12043 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__dfrtn_1_2/a_543_47# 0.00fF
C12044 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# 0.00fF
C12045 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__or3_1_0/C 0.01fF
C12046 sky130_fd_sc_hd__inv_1_12/A sky130_fd_sc_hd__inv_1_8/A 0.01fF
C12047 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__inv_1_39/A 0.01fF
C12048 sky130_fd_sc_hd__dfrtn_1_34/a_1217_47# DONE 0.00fF
C12049 sky130_fd_sc_hd__inv_1_41/Y SEL_CONV_TIME[3] 0.21fF
C12050 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_24/a_543_47# -0.00fF
C12051 sky130_fd_sc_hd__dfrtn_1_27/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12052 DOUT[9] sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C12053 sky130_fd_sc_hd__dfrtn_1_38/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12054 sky130_fd_sc_hd__dfrtp_1_3/a_651_413# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C12055 sky130_fd_sc_hd__inv_1_1/A DOUT[22] 0.00fF
C12056 sky130_fd_sc_hd__inv_1_22/Y DOUT[12] 0.00fF
C12057 sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C12058 DOUT[1] sky130_fd_sc_hd__dfrtn_1_22/a_448_47# 0.00fF
C12059 sky130_fd_sc_hd__inv_1_6/A VIN 0.16fF
C12060 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C12061 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# DOUT[21] 0.00fF
C12062 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_41/a_761_289# 0.03fF
C12063 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_0/Y 0.03fF
C12064 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# DOUT[23] 0.00fF
C12065 sky130_fd_sc_hd__inv_1_52/A DOUT[4] 0.02fF
C12066 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C12067 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# DOUT[14] 0.00fF
C12068 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# DOUT[19] 0.02fF
C12069 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C12070 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# 0.01fF
C12071 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_15/a_761_289# 0.00fF
C12072 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C12073 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C12074 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_448_47# 0.00fF
C12075 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C12076 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C12077 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C12078 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# sky130_fd_sc_hd__inv_1_42/Y 0.02fF
C12079 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C12080 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# sky130_fd_sc_hd__nor3_1_0/a_109_297# 0.00fF
C12081 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C12082 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__inv_1_54/Y 0.00fF
C12083 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C12084 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C12085 sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# VDD 0.07fF
C12086 sky130_fd_sc_hd__dfrtn_1_36/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12087 sky130_fd_sc_hd__inv_1_41/Y SEL_CONV_TIME[2] 0.37fF
C12088 sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C12089 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# 0.00fF
C12090 sky130_fd_sc_hd__dfrtn_1_12/a_761_289# sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# 0.00fF
C12091 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__dfrtn_1_13/a_27_47# 0.00fF
C12092 sky130_fd_sc_hd__dfrtn_1_0/a_639_47# DOUT[18] 0.00fF
C12093 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__or2b_1_0/X 0.02fF
C12094 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# SEL_CONV_TIME[3] 0.00fF
C12095 sky130_fd_sc_hd__nor3_2_3/a_27_297# sky130_fd_sc_hd__dfrtn_1_42/a_27_47# 0.00fF
C12096 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# 0.01fF
C12097 sky130_fd_sc_hd__dfrtn_1_26/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12098 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_13/a_27_47# 0.00fF
C12099 sky130_fd_sc_hd__dfrtn_1_0/a_651_413# sky130_fd_sc_hd__nor3_1_0/A 0.01fF
C12100 sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C12101 sky130_fd_sc_hd__dfrtn_1_34/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12102 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_27/a_639_47# 0.00fF
C12103 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__o2111a_2_0/X 0.01fF
C12104 sky130_fd_sc_hd__nand3b_1_1/Y sky130_fd_sc_hd__inv_1_44/A 0.12fF
C12105 sky130_fd_sc_hd__nor3_1_19/Y SEL_CONV_TIME[1] 0.30fF
C12106 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C12107 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_1/a_805_47# 0.00fF
C12108 sky130_fd_sc_hd__dfrtn_1_28/a_448_47# RESET_COUNTERn 0.00fF
C12109 sky130_fd_sc_hd__dfrtn_1_28/a_1217_47# DOUT[21] 0.00fF
C12110 sky130_fd_sc_hd__dfrtn_1_39/a_651_413# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C12111 sky130_fd_sc_hd__dfrtn_1_30/a_651_413# sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C12112 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__nand2_1_1/Y 0.01fF
C12113 sky130_fd_sc_hd__mux4_1_0/a_668_97# SEL_CONV_TIME[0] 0.00fF
C12114 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# 0.00fF
C12115 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12116 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# DOUT[21] 0.01fF
C12117 sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# VDD 0.07fF
C12118 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C12119 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_12/a_193_47# 0.00fF
C12120 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# sky130_fd_sc_hd__inv_1_39/A 0.02fF
C12121 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C12122 DOUT[4] sky130_fd_sc_hd__dfrtn_1_24/a_27_47# 0.00fF
C12123 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_761_289# 0.00fF
C12124 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_193_47# 0.00fF
C12125 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# SEL_CONV_TIME[2] 0.03fF
C12126 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# VIN 0.00fF
C12127 sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# 0.00fF
C12128 sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.00fF
C12129 sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# DOUT[22] 0.00fF
C12130 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C12131 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_448_47# 0.00fF
C12132 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C12133 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C12134 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C12135 sky130_fd_sc_hd__inv_1_7/A RESET_COUNTERn 0.63fF
C12136 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C12137 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C12138 sky130_fd_sc_hd__inv_1_31/A DOUT[2] 0.01fF
C12139 sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# sky130_fd_sc_hd__inv_1_9/A 0.00fF
C12140 sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# RESET_COUNTERn 0.01fF
C12141 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# SEL_CONV_TIME[0] 0.00fF
C12142 sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# DOUT[2] 0.01fF
C12143 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__inv_1_29/Y 0.00fF
C12144 DOUT[1] sky130_fd_sc_hd__dfrtn_1_23/a_651_413# 0.00fF
C12145 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_761_289# 0.00fF
C12146 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.00fF
C12147 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C12148 sky130_fd_sc_hd__or2_2_0/X DOUT[0] 0.00fF
C12149 sky130_fd_sc_hd__dfrtn_1_32/a_193_47# VDD 0.09fF
C12150 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_25/a_805_47# 0.00fF
C12151 sky130_fd_sc_hd__dfrtn_1_22/a_1217_47# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C12152 sky130_fd_sc_hd__inv_1_44/A sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C12153 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# -0.00fF
C12154 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# -0.00fF
C12155 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# -0.00fF
C12156 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C12157 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_38/a_761_289# 0.00fF
C12158 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C12159 sky130_fd_sc_hd__dfrtn_1_31/a_1270_413# SEL_CONV_TIME[1] 0.00fF
C12160 sky130_fd_sc_hd__mux4_1_0/a_757_363# RESET_COUNTERn 0.01fF
C12161 VIN out 0.83fF
C12162 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.01fF
C12163 sky130_fd_sc_hd__dfrtn_1_10/a_639_47# RESET_COUNTERn 0.00fF
C12164 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C12165 CLK_REF sky130_fd_sc_hd__nor3_2_3/B 0.24fF
C12166 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_24/a_27_47# 0.01fF
C12167 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_19/a_805_47# 0.00fF
C12168 sky130_fd_sc_hd__or3b_2_0/a_472_297# sky130_fd_sc_hd__dfrtn_1_31/a_543_47# 0.00fF
C12169 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_31/a_448_47# 0.00fF
C12170 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_1108_47# 0.00fF
C12171 sky130_fd_sc_hd__dfrtn_1_21/a_761_289# sky130_fd_sc_hd__inv_1_35/A 0.01fF
C12172 sky130_fd_sc_hd__inv_1_52/A outb 0.02fF
C12173 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# DOUT[19] 0.00fF
C12174 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__inv_1_48/A 0.01fF
C12175 sky130_fd_sc_hd__nor3_1_14/a_109_297# outb 0.00fF
C12176 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__dfrtn_1_15/a_805_47# 0.00fF
C12177 sky130_fd_sc_hd__dfrtn_1_17/a_639_47# VDD 0.00fF
C12178 sky130_fd_sc_hd__dfrtn_1_28/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C12179 sky130_fd_sc_hd__dfrtn_1_17/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12180 sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C12181 sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12182 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__nor3_1_0/a_193_297# 0.00fF
C12183 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# sky130_fd_sc_hd__nor3_1_0/a_109_297# 0.00fF
C12184 sky130_fd_sc_hd__dfrtn_1_32/a_27_47# sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# -0.00fF
C12185 sky130_fd_sc_hd__dfrtn_1_32/a_761_289# sky130_fd_sc_hd__dfrtn_1_32/a_543_47# -0.00fF
C12186 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# 0.00fF
C12187 DOUT[2] sky130_fd_sc_hd__inv_1_33/A 0.43fF
C12188 sky130_fd_sc_hd__nor3_2_3/a_281_297# sky130_fd_sc_hd__dfrtn_1_42/a_805_47# 0.00fF
C12189 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# 0.00fF
C12190 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C12191 sky130_fd_sc_hd__dfrtn_1_22/a_1108_47# sky130_fd_sc_hd__inv_1_37/A 0.01fF
C12192 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__dfrtn_1_31/a_27_47# 0.00fF
C12193 sky130_fd_sc_hd__inv_1_53/Y RESET_COUNTERn 0.18fF
C12194 DOUT[17] DOUT[18] 0.33fF
C12195 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__dfrtn_1_19/a_448_47# 0.00fF
C12196 sky130_fd_sc_hd__dfrtn_1_3/a_639_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C12197 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__dfrtn_1_30/a_761_289# -0.00fF
C12198 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.00fF
C12199 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C12200 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C12201 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C12202 sky130_fd_sc_hd__nor3_1_11/a_193_297# sky130_fd_sc_hd__dfrtn_1_7/a_193_47# 0.00fF
C12203 sky130_fd_sc_hd__inv_1_9/Y sky130_fd_sc_hd__inv_1_9/A 0.00fF
C12204 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfrtn_1_41/a_761_289# 0.00fF
C12205 sky130_fd_sc_hd__dfrtn_1_31/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12206 sky130_fd_sc_hd__dfrtn_1_31/a_651_413# VDD 0.01fF
C12207 sky130_fd_sc_hd__dfrtn_1_3/a_761_289# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C12208 sky130_fd_sc_hd__mux4_2_0/a_1279_413# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C12209 sky130_fd_sc_hd__nand3b_1_0/Y VDD 0.31fF
C12210 sky130_fd_sc_hd__dfrtn_1_38/a_761_289# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C12211 sky130_fd_sc_hd__dfrtn_1_28/a_761_289# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C12212 sky130_fd_sc_hd__mux4_2_0/a_872_316# SEL_CONV_TIME[0] 0.02fF
C12213 sky130_fd_sc_hd__dfrtn_1_0/a_805_47# RESET_COUNTERn 0.00fF
C12214 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C12215 sky130_fd_sc_hd__dfrtn_1_35/a_448_47# RESET_COUNTERn 0.00fF
C12216 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_448_47# -0.00fF
C12217 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# sky130_fd_sc_hd__dfrtn_1_31/a_1108_47# -0.00fF
C12218 sky130_fd_sc_hd__dfrtn_1_29/a_639_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C12219 sky130_fd_sc_hd__dfrtn_1_23/a_1462_47# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C12220 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C12221 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# DOUT[3] 0.00fF
C12222 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_1462_47# 0.00fF
C12223 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# 0.00fF
C12224 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_30/a_805_47# 0.00fF
C12225 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# RESET_COUNTERn 0.00fF
C12226 sky130_fd_sc_hd__dfrtp_1_3/a_761_289# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C12227 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C12228 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_761_289# 0.00fF
C12229 sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C12230 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_19/a_639_47# 0.00fF
C12231 sky130_fd_sc_hd__dfrtn_1_40/a_1270_413# sky130_fd_sc_hd__inv_1_31/A 0.00fF
C12232 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__inv_1_43/Y 0.01fF
C12233 sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# SEL_CONV_TIME[0] 0.00fF
C12234 sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C12235 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_38/a_639_47# 0.00fF
C12236 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C12237 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_18/a_805_47# 0.00fF
C12238 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_40/a_27_47# 0.00fF
C12239 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_18/a_1217_47# 0.00fF
C12240 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_18/a_651_413# 0.00fF
C12241 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_1462_47# 0.00fF
C12242 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C12243 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C12244 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# RESET_COUNTERn 0.03fF
C12245 sky130_fd_sc_hd__dfrtn_1_32/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12246 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C12247 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__dfrtn_1_29/a_761_289# 0.00fF
C12248 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C12249 sky130_fd_sc_hd__dfrtn_1_32/a_1462_47# VDD 0.00fF
C12250 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12251 sky130_fd_sc_hd__dfrtn_1_7/a_651_413# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C12252 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# VDD 0.11fF
C12253 sky130_fd_sc_hd__dfrtn_1_3/a_805_47# DOUT[11] 0.00fF
C12254 sky130_fd_sc_hd__dfrtn_1_4/a_805_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C12255 sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C12256 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__dfrtn_1_1/a_543_47# -0.00fF
C12257 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# -0.00fF
C12258 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# SEL_CONV_TIME[1] 0.00fF
C12259 sky130_fd_sc_hd__dfrtn_1_36/a_805_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C12260 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__inv_1_7/A 0.28fF
C12261 sky130_fd_sc_hd__o311a_1_0/a_81_21# RESET_COUNTERn 0.00fF
C12262 sky130_fd_sc_hd__dfrtp_1_3/a_1270_413# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C12263 sky130_fd_sc_hd__inv_1_6/Y RESET_COUNTERn 0.04fF
C12264 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C12265 sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# SEL_CONV_TIME[0] 0.00fF
C12266 sky130_fd_sc_hd__or2b_1_0/a_301_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12267 sky130_fd_sc_hd__mux4_2_0/a_193_369# RESET_COUNTERn 0.00fF
C12268 sky130_fd_sc_hd__or3_1_0/X sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C12269 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__nor3_2_3/C 0.13fF
C12270 sky130_fd_sc_hd__dfrtn_1_23/a_448_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C12271 sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# sky130_fd_sc_hd__dfrtn_1_28/a_448_47# 0.00fF
C12272 sky130_fd_sc_hd__nor3_1_18/a_109_297# sky130_fd_sc_hd__nor3_2_2/a_27_297# 0.00fF
C12273 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# 0.01fF
C12274 sky130_fd_sc_hd__nor3_1_15/a_109_297# sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.00fF
C12275 sky130_fd_sc_hd__inv_1_14/A sky130_fd_sc_hd__inv_1_8/A 0.01fF
C12276 sky130_fd_sc_hd__nor3_1_4/A DOUT[7] 0.23fF
C12277 sky130_fd_sc_hd__nor3_1_15/a_109_297# sky130_fd_sc_hd__inv_1_9/A 0.00fF
C12278 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C12279 sky130_fd_sc_hd__dfrtn_1_42/a_1270_413# sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C12280 sky130_fd_sc_hd__dfrtn_1_4/a_448_47# DOUT[11] 0.00fF
C12281 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# RESET_COUNTERn 0.05fF
C12282 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__dfrtn_1_33/a_543_47# -0.00fF
C12283 sky130_fd_sc_hd__dfrtn_1_0/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12284 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12285 sky130_fd_sc_hd__inv_1_45/Y RESET_COUNTERn 0.21fF
C12286 sky130_fd_sc_hd__dfrtn_1_35/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C12287 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# VDD 0.00fF
C12288 sky130_fd_sc_hd__dfrtn_1_40/a_1270_413# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C12289 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# RESET_COUNTERn 0.03fF
C12290 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_34/a_448_47# 0.00fF
C12291 sky130_fd_sc_hd__inv_1_11/Y sky130_fd_sc_hd__inv_1_5/A 0.00fF
C12292 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__nor3_2_1/a_27_297# 0.00fF
C12293 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.62fF
C12294 DOUT[4] sky130_fd_sc_hd__dfrtn_1_30/a_805_47# 0.00fF
C12295 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# VDD 0.06fF
C12296 sky130_fd_sc_hd__nand3b_1_0/a_316_47# RESET_COUNTERn 0.00fF
C12297 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__or2_2_0/X 0.01fF
C12298 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__dfrtn_1_5/a_639_47# 0.00fF
C12299 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C12300 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C12301 DOUT[13] sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C12302 sky130_fd_sc_hd__dfrtn_1_19/a_651_413# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C12303 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__inv_1_8/Y 0.01fF
C12304 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.00fF
C12305 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__o211a_1_1/a_215_47# 0.00fF
C12306 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__o211a_1_1/a_297_297# 0.00fF
C12307 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.00fF
C12308 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C12309 sky130_fd_sc_hd__dfrtn_1_25/a_805_47# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C12310 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__o211a_1_1/X 0.00fF
C12311 sky130_fd_sc_hd__inv_1_15/A DOUT[7] 0.00fF
C12312 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C12313 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C12314 sky130_fd_sc_hd__dfrtn_1_27/a_543_47# DOUT[21] 0.00fF
C12315 sky130_fd_sc_hd__nor3_1_4/A sky130_fd_sc_hd__inv_1_12/A 0.04fF
C12316 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__inv_1_13/A 0.01fF
C12317 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C12318 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_1/a_448_47# 0.00fF
C12319 sky130_fd_sc_hd__dfrtn_1_11/a_761_289# sky130_fd_sc_hd__inv_1_12/A 0.01fF
C12320 sky130_fd_sc_hd__o211a_1_0/a_297_297# DOUT[23] 0.00fF
C12321 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__nor3_1_2/a_109_297# 0.00fF
C12322 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_25/a_543_47# 0.00fF
C12323 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__dfrtn_1_25/a_761_289# 0.00fF
C12324 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__dfrtn_1_25/a_193_47# 0.00fF
C12325 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_25/a_448_47# 0.00fF
C12326 sky130_fd_sc_hd__dfrtp_1_3/a_448_47# sky130_fd_sc_hd__dfrtn_1_17/a_651_413# 0.00fF
C12327 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_1462_47# 0.00fF
C12328 sky130_fd_sc_hd__dfrtp_1_3/a_761_289# sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# 0.00fF
C12329 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_32/a_193_47# 0.00fF
C12330 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C12331 sky130_fd_sc_hd__nor3_2_0/A DOUT[22] 0.00fF
C12332 sky130_fd_sc_hd__nor3_1_15/a_109_297# sky130_fd_sc_hd__dfrtn_1_32/a_27_47# 0.00fF
C12333 sky130_fd_sc_hd__dfrtn_1_12/a_639_47# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C12334 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C12335 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C12336 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.00fF
C12337 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# sky130_fd_sc_hd__mux4_2_0/a_193_369# 0.00fF
C12338 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtp_1_2/a_651_413# -0.00fF
C12339 sky130_fd_sc_hd__dfrtn_1_4/a_761_289# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C12340 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C12341 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__dfrtn_1_29/a_805_47# 0.00fF
C12342 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C12343 sky130_fd_sc_hd__dfrtn_1_4/a_639_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C12344 DOUT[22] DOUT[17] 0.03fF
C12345 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__nand3b_1_1/Y 0.01fF
C12346 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# 0.00fF
C12347 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C12348 sky130_fd_sc_hd__o2111a_2_0/a_386_47# sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# 0.00fF
C12349 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__dfrtn_1_24/a_761_289# 0.00fF
C12350 CLK_REF DOUT[0] 0.00fF
C12351 sky130_fd_sc_hd__dfrtp_1_3/a_1462_47# VDD 0.00fF
C12352 sky130_fd_sc_hd__dfrtp_1_3/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12353 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# RESET_COUNTERn 0.05fF
C12354 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# sky130_fd_sc_hd__dfrtn_1_26/a_761_289# 0.00fF
C12355 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_543_47# 0.00fF
C12356 sky130_fd_sc_hd__nor3_1_18/a_193_297# DOUT[15] 0.00fF
C12357 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C12358 sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# sky130_fd_sc_hd__or3b_2_0/X 0.01fF
C12359 sky130_fd_sc_hd__dfrtn_1_22/a_543_47# VDD 0.06fF
C12360 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12361 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# RESET_COUNTERn 0.33fF
C12362 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# 0.01fF
C12363 DOUT[1] sky130_fd_sc_hd__dfrtn_1_42/a_193_47# 0.00fF
C12364 sky130_fd_sc_hd__inv_1_53/A sky130_fd_sc_hd__inv_1_41/Y 0.02fF
C12365 SEL_CONV_TIME[0] SEL_CONV_TIME[1] 2.27fF
C12366 sky130_fd_sc_hd__inv_1_53/Y SEL_CONV_TIME[2] 0.00fF
C12367 sky130_fd_sc_hd__nor3_1_5/A DOUT[21] 0.01fF
C12368 sky130_fd_sc_hd__dfrtn_1_28/a_1108_47# sky130_fd_sc_hd__inv_1_48/A 0.01fF
C12369 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C12370 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# 0.00fF
C12371 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C12372 DOUT[4] sky130_fd_sc_hd__dfrtn_1_34/a_448_47# 0.00fF
C12373 sky130_fd_sc_hd__or3_1_0/C RESET_COUNTERn 0.25fF
C12374 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C12375 sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# 0.00fF
C12376 sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# 0.00fF
C12377 sky130_fd_sc_hd__nor3_1_3/a_193_297# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C12378 sky130_fd_sc_hd__nor3_1_2/a_109_297# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C12379 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__dfrtn_1_6/a_27_47# 0.00fF
C12380 DOUT[1] sky130_fd_sc_hd__inv_1_38/A 0.00fF
C12381 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# sky130_fd_sc_hd__inv_1_40/A 0.03fF
C12382 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C12383 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C12384 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_805_47# -0.00fF
C12385 sky130_fd_sc_hd__or2b_1_0/X RESET_COUNTERn 0.11fF
C12386 sky130_fd_sc_hd__dfrtn_1_11/a_1217_47# RESET_COUNTERn 0.00fF
C12387 sky130_fd_sc_hd__o311a_1_0/a_81_21# SEL_CONV_TIME[3] 0.02fF
C12388 sky130_fd_sc_hd__dfrtn_1_8/a_193_47# sky130_fd_sc_hd__inv_1_9/A 0.00fF
C12389 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__inv_1_6/Y 0.01fF
C12390 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_10/a_448_47# 0.00fF
C12391 sky130_fd_sc_hd__dfrtp_1_1/a_448_47# DOUT[23] 0.00fF
C12392 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C12393 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C12394 sky130_fd_sc_hd__nor3_1_0/a_109_297# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C12395 sky130_fd_sc_hd__dfrtn_1_8/a_448_47# DOUT[12] 0.00fF
C12396 sky130_fd_sc_hd__mux4_2_0/a_193_369# SEL_CONV_TIME[3] 0.00fF
C12397 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__nor3_2_0/A 0.01fF
C12398 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C12399 sky130_fd_sc_hd__dfrtn_1_16/a_193_47# VDD 0.08fF
C12400 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C12401 sky130_fd_sc_hd__o211a_1_0/a_79_21# sky130_fd_sc_hd__inv_1_26/A 0.00fF
C12402 sky130_fd_sc_hd__nor3_1_6/a_193_297# VDD 0.00fF
C12403 sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12404 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__inv_1_53/A 0.02fF
C12405 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__dfrtp_1_3/a_1108_47# -0.00fF
C12406 sky130_fd_sc_hd__dfrtp_1_3/a_761_289# sky130_fd_sc_hd__dfrtp_1_3/a_543_47# -0.00fF
C12407 sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12408 CLK_REF sky130_fd_sc_hd__dfrtn_1_19/a_448_47# 0.00fF
C12409 sky130_fd_sc_hd__nor3_2_2/a_27_297# VDD 0.06fF
C12410 sky130_fd_sc_hd__nor3_1_3/a_193_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12411 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# sky130_fd_sc_hd__inv_1_1/A 0.01fF
C12412 sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# sky130_fd_sc_hd__dfrtn_1_18/a_651_413# 0.00fF
C12413 sky130_fd_sc_hd__dfrtn_1_20/a_1462_47# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C12414 sky130_fd_sc_hd__dfrtn_1_20/a_1217_47# sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.00fF
C12415 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C12416 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# 0.00fF
C12417 sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C12418 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__nand3b_1_0/a_53_93# 0.00fF
C12419 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# sky130_fd_sc_hd__inv_1_3/A 0.02fF
C12420 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# DOUT[2] 0.00fF
C12421 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C12422 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_34/a_448_47# 0.00fF
C12423 sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C12424 sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# sky130_fd_sc_hd__dfrtn_1_36/a_651_413# 0.00fF
C12425 sky130_fd_sc_hd__dfrtn_1_23/a_1462_47# sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C12426 sky130_fd_sc_hd__dfrtn_1_23/a_1217_47# sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C12427 sky130_fd_sc_hd__dfrtn_1_21/a_543_47# DOUT[2] 0.00fF
C12428 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_543_47# -0.00fF
C12429 sky130_fd_sc_hd__dfrtn_1_27/a_639_47# RESET_COUNTERn 0.00fF
C12430 sky130_fd_sc_hd__dfrtn_1_38/a_805_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C12431 sky130_fd_sc_hd__o311a_1_0/a_81_21# SEL_CONV_TIME[2] 0.01fF
C12432 sky130_fd_sc_hd__inv_1_43/A sky130_fd_sc_hd__nor3_2_3/B 0.08fF
C12433 sky130_fd_sc_hd__dfrtn_1_35/a_805_47# sky130_fd_sc_hd__inv_1_38/A 0.00fF
C12434 DOUT[13] sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C12435 sky130_fd_sc_hd__nand3b_1_0/a_316_47# SEL_CONV_TIME[3] 0.00fF
C12436 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C12437 sky130_fd_sc_hd__mux4_2_0/a_193_369# SEL_CONV_TIME[2] 0.00fF
C12438 sky130_fd_sc_hd__nor3_1_11/a_109_297# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C12439 sky130_fd_sc_hd__nor3_1_11/a_193_297# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C12440 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# VDD 0.09fF
C12441 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_32/a_1462_47# 0.00fF
C12442 sky130_fd_sc_hd__dfrtn_1_30/a_651_413# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C12443 sky130_fd_sc_hd__nor3_2_0/a_281_297# sky130_fd_sc_hd__dfrtn_1_12/a_448_47# 0.00fF
C12444 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# -0.00fF
C12445 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# -0.00fF
C12446 DOUT[13] sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# 0.01fF
C12447 sky130_fd_sc_hd__dfrtn_1_38/a_1270_413# DOUT[2] 0.00fF
C12448 sky130_fd_sc_hd__dfrtn_1_37/a_1270_413# sky130_fd_sc_hd__mux4_2_0/a_872_316# 0.00fF
C12449 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# sky130_fd_sc_hd__mux4_2_0/a_1064_47# 0.00fF
C12450 sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C12451 sky130_fd_sc_hd__dfrtn_1_37/a_805_47# sky130_fd_sc_hd__mux4_2_0/a_600_345# 0.00fF
C12452 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C12453 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C12454 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# sky130_fd_sc_hd__mux4_2_0/a_397_47# 0.00fF
C12455 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_38/a_761_289# 0.00fF
C12456 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__nor3_2_0/a_281_297# 0.00fF
C12457 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# VDD 0.18fF
C12458 sky130_fd_sc_hd__mux4_2_0/a_397_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12459 DOUT[16] RESET_COUNTERn 0.01fF
C12460 sky130_fd_sc_hd__dfrtn_1_36/a_193_47# RESET_COUNTERn 0.31fF
C12461 sky130_fd_sc_hd__dfrtn_1_36/a_448_47# DOUT[21] 0.00fF
C12462 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# sky130_fd_sc_hd__inv_1_32/A 0.01fF
C12463 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# sky130_fd_sc_hd__or2_2_0/B 0.01fF
C12464 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# RESET_COUNTERn 0.00fF
C12465 sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C12466 sky130_fd_sc_hd__dfrtn_1_14/a_448_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C12467 sky130_fd_sc_hd__dfrtn_1_33/a_639_47# sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# 0.00fF
C12468 sky130_fd_sc_hd__dfrtn_1_33/a_805_47# sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# 0.00fF
C12469 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# VDD 0.01fF
C12470 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12471 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# 0.00fF
C12472 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# 0.00fF
C12473 sky130_fd_sc_hd__dfrtn_1_22/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12474 sky130_fd_sc_hd__nor3_1_12/a_109_297# sky130_fd_sc_hd__dfrtn_1_8/a_448_47# 0.00fF
C12475 sky130_fd_sc_hd__nor3_1_12/a_193_297# sky130_fd_sc_hd__dfrtn_1_8/a_1108_47# 0.00fF
C12476 sky130_fd_sc_hd__dfrtn_1_11/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12477 sky130_fd_sc_hd__dfrtn_1_12/a_1462_47# RESET_COUNTERn 0.00fF
C12478 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_805_47# -0.00fF
C12479 sky130_fd_sc_hd__dfrtn_1_20/a_543_47# sky130_fd_sc_hd__dfrtn_1_21/a_1462_47# 0.00fF
C12480 DOUT[1] sky130_fd_sc_hd__dfrtn_1_42/a_1462_47# 0.00fF
C12481 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C12482 sky130_fd_sc_hd__nor3_1_15/a_193_297# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C12483 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C12484 sky130_fd_sc_hd__inv_1_30/Y sky130_fd_sc_hd__inv_1_33/A 0.00fF
C12485 sky130_fd_sc_hd__inv_1_35/Y DOUT[2] 0.00fF
C12486 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__dfrtn_1_25/a_448_47# 0.00fF
C12487 sky130_fd_sc_hd__or2_2_0/A RESET_COUNTERn 0.28fF
C12488 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C12489 sky130_fd_sc_hd__dfrtn_1_18/a_1270_413# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C12490 sky130_fd_sc_hd__nor3_1_7/a_193_297# DOUT[6] 0.00fF
C12491 sky130_fd_sc_hd__nor3_1_7/a_109_297# DOUT[7] 0.00fF
C12492 sky130_fd_sc_hd__dfrtn_1_27/a_193_47# DOUT[23] 0.00fF
C12493 sky130_fd_sc_hd__dfrtp_1_0/a_639_47# sky130_fd_sc_hd__dfrtp_1_1/a_193_47# 0.00fF
C12494 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__dfrtp_1_1/a_805_47# 0.00fF
C12495 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/a_639_47# 0.00fF
C12496 sky130_fd_sc_hd__inv_1_32/A sky130_fd_sc_hd__inv_1_32/Y 0.02fF
C12497 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# DOUT[0] 0.00fF
C12498 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# 0.00fF
C12499 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.00fF
C12500 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_761_289# 0.00fF
C12501 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.01fF
C12502 sky130_fd_sc_hd__dfrtn_1_0/a_1462_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C12503 sky130_fd_sc_hd__dfrtn_1_8/a_1462_47# sky130_fd_sc_hd__inv_1_9/A 0.00fF
C12504 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__dfrtn_1_13/a_761_289# 0.00fF
C12505 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__dfrtn_1_13/a_193_47# 0.00fF
C12506 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__inv_1_47/Y 0.00fF
C12507 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# sky130_fd_sc_hd__nor3_1_4/a_193_297# 0.00fF
C12508 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__nor3_1_4/a_109_297# 0.00fF
C12509 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C12510 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_20/a_27_47# 0.01fF
C12511 sky130_fd_sc_hd__or3_1_0/C SEL_CONV_TIME[3] 0.01fF
C12512 sky130_fd_sc_hd__dfrtn_1_26/a_651_413# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C12513 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C12514 sky130_fd_sc_hd__dfrtn_1_5/a_805_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C12515 sky130_fd_sc_hd__mux4_2_0/a_1281_47# SEL_CONV_TIME[3] 0.00fF
C12516 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# DOUT[11] 0.00fF
C12517 sky130_fd_sc_hd__dfrtn_1_16/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12518 sky130_fd_sc_hd__dfrtn_1_27/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12519 sky130_fd_sc_hd__dfrtn_1_16/a_1462_47# VDD 0.00fF
C12520 sky130_fd_sc_hd__dfrtn_1_8/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C12521 sky130_fd_sc_hd__dfrtn_1_8/a_1270_413# VDD 0.00fF
C12522 sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C12523 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__nor3_1_19/a_109_297# 0.00fF
C12524 sky130_fd_sc_hd__dfrtn_1_34/a_543_47# sky130_fd_sc_hd__inv_1_49/A 0.02fF
C12525 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__dfrtn_1_29/a_448_47# -0.00fF
C12526 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_651_413# -0.00fF
C12527 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__inv_1_7/A 0.01fF
C12528 DOUT[13] sky130_fd_sc_hd__dfrtn_1_34/a_193_47# 0.00fF
C12529 sky130_fd_sc_hd__dfrtn_1_24/a_651_413# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C12530 sky130_fd_sc_hd__dfrtn_1_32/a_761_289# DOUT[21] 0.00fF
C12531 sky130_fd_sc_hd__nor3_1_19/Y DOUT[21] 0.01fF
C12532 sky130_fd_sc_hd__or2b_1_0/X SEL_CONV_TIME[3] 0.00fF
C12533 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C12534 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__dfrtn_1_34/a_27_47# 0.00fF
C12535 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_20/a_805_47# 0.00fF
C12536 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# CLK_REF 0.02fF
C12537 sky130_fd_sc_hd__dfrtn_1_19/a_27_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C12538 DOUT[4] sky130_fd_sc_hd__dfrtn_1_10/a_761_289# 0.00fF
C12539 sky130_fd_sc_hd__dfrtn_1_31/a_639_47# SEL_CONV_TIME[0] 0.00fF
C12540 sky130_fd_sc_hd__dfrtn_1_25/a_448_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C12541 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C12542 sky130_fd_sc_hd__or3b_2_0/a_472_297# RESET_COUNTERn 0.00fF
C12543 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12544 sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C12545 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__inv_1_44/A 0.01fF
C12546 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# DOUT[14] 0.00fF
C12547 DOUT[12] sky130_fd_sc_hd__nor3_2_3/B 1.27fF
C12548 sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# sky130_fd_sc_hd__or3_1_0/C 0.01fF
C12549 sky130_fd_sc_hd__dfrtn_1_12/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12550 sky130_fd_sc_hd__or3_1_0/a_183_297# sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# 0.00fF
C12551 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C12552 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__inv_1_32/A 0.01fF
C12553 sky130_fd_sc_hd__nor3_2_1/a_27_297# DOUT[15] 0.00fF
C12554 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_3/a_1270_413# 0.00fF
C12555 sky130_fd_sc_hd__dfrtn_1_7/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12556 sky130_fd_sc_hd__dfrtn_1_7/a_1217_47# VDD 0.00fF
C12557 sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# RESET_COUNTERn 0.02fF
C12558 sky130_fd_sc_hd__nor3_1_19/Y sky130_fd_sc_hd__o311a_1_0/A3 0.01fF
C12559 sky130_fd_sc_hd__or2b_1_0/X SEL_CONV_TIME[2] 0.00fF
C12560 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# DOUT[14] 0.00fF
C12561 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__inv_1_54/A 0.03fF
C12562 sky130_fd_sc_hd__dfrtn_1_9/a_651_413# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C12563 sky130_fd_sc_hd__dfrtn_1_36/a_1462_47# RESET_COUNTERn 0.00fF
C12564 sky130_fd_sc_hd__dfrtn_1_3/a_805_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C12565 CLK_REF DOUT[2] 0.02fF
C12566 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_1283_21# 0.02fF
C12567 sky130_fd_sc_hd__dfrtn_1_21/a_448_47# sky130_fd_sc_hd__dfrtn_1_19/a_1108_47# 0.00fF
C12568 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__inv_1_7/A 0.01fF
C12569 sky130_fd_sc_hd__nand3b_1_0/a_232_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C12570 sky130_fd_sc_hd__nor3_1_1/a_193_297# VDD 0.00fF
C12571 sky130_fd_sc_hd__dfrtn_1_0/a_543_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C12572 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.00fF
C12573 sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# sky130_fd_sc_hd__inv_1_11/Y 0.03fF
C12574 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# 0.00fF
C12575 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C12576 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# 0.00fF
C12577 sky130_fd_sc_hd__nor3_2_3/C lc_out 0.11fF
C12578 sky130_fd_sc_hd__dfrtn_1_31/a_543_47# RESET_COUNTERn 0.01fF
C12579 sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# sky130_fd_sc_hd__inv_1_53/A 0.01fF
C12580 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C12581 sky130_fd_sc_hd__dfrtn_1_9/a_543_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C12582 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12583 sky130_fd_sc_hd__or2_2_0/a_39_297# sky130_fd_sc_hd__dfrtn_1_19/a_543_47# 0.00fF
C12584 sky130_fd_sc_hd__dfrtn_1_27/a_1462_47# DOUT[23] 0.00fF
C12585 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C12586 DONE sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C12587 sky130_fd_sc_hd__dfrtn_1_4/a_448_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C12588 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C12589 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C12590 sky130_fd_sc_hd__dfrtn_1_25/a_448_47# sky130_fd_sc_hd__dfrtn_1_27/a_651_413# 0.00fF
C12591 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_1462_47# 0.00fF
C12592 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# sky130_fd_sc_hd__dfrtn_1_27/a_1217_47# 0.00fF
C12593 sky130_fd_sc_hd__dfrtn_1_20/a_761_289# DOUT[2] 0.01fF
C12594 sky130_fd_sc_hd__o311a_1_0/a_266_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C12595 sky130_fd_sc_hd__inv_1_14/A sky130_fd_sc_hd__inv_1_15/A 0.00fF
C12596 sky130_fd_sc_hd__dfrtn_1_42/a_1217_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C12597 sky130_fd_sc_hd__inv_1_24/A VIN 0.13fF
C12598 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__inv_1_3/A 0.76fF
C12599 sky130_fd_sc_hd__nor3_1_10/a_193_297# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C12600 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# DONE 0.00fF
C12601 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__inv_1_33/A 0.01fF
C12602 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__inv_1_37/A 0.02fF
C12603 sky130_fd_sc_hd__dfrtn_1_19/a_1108_47# sky130_fd_sc_hd__inv_1_35/A 0.00fF
C12604 sky130_fd_sc_hd__inv_1_45/A RESET_COUNTERn 0.23fF
C12605 sky130_fd_sc_hd__nor3_1_12/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12606 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12607 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# 0.01fF
C12608 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C12609 sky130_fd_sc_hd__inv_1_33/Y RESET_COUNTERn 0.01fF
C12610 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C12611 DOUT[13] sky130_fd_sc_hd__dfrtn_1_34/a_1462_47# 0.00fF
C12612 sky130_fd_sc_hd__dfrtn_1_32/a_1270_413# RESET_COUNTERn 0.00fF
C12613 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# SEL_CONV_TIME[0] 0.02fF
C12614 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__dfrtn_1_33/a_761_289# 0.00fF
C12615 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__dfrtn_1_33/a_27_47# 0.00fF
C12616 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_33/a_193_47# 0.00fF
C12617 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# 0.00fF
C12618 sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__dfrtn_1_33/a_543_47# 0.00fF
C12619 sky130_fd_sc_hd__o311a_1_0/a_81_21# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C12620 DOUT[4] DOUT[1] 0.03fF
C12621 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# -0.00fF
C12622 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# -0.00fF
C12623 sky130_fd_sc_hd__dfrtn_1_8/a_651_413# sky130_fd_sc_hd__inv_1_9/Y 0.00fF
C12624 sky130_fd_sc_hd__dfrtn_1_21/a_1462_47# sky130_fd_sc_hd__inv_1_35/A 0.00fF
C12625 sky130_fd_sc_hd__dfrtn_1_28/a_448_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C12626 sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# CLK_REF 0.00fF
C12627 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__inv_1_13/A 0.01fF
C12628 sky130_fd_sc_hd__dfrtn_1_17/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12629 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# outb 0.00fF
C12630 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__dfrtn_1_22/a_639_47# -0.00fF
C12631 sky130_fd_sc_hd__dfrtn_1_36/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12632 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# 0.00fF
C12633 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C12634 sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C12635 sky130_fd_sc_hd__or2b_1_0/a_219_297# RESET_COUNTERn 0.00fF
C12636 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C12637 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# VDD 0.01fF
C12638 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_4/Y 0.01fF
C12639 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_8/A 0.00fF
C12640 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__nor3_2_3/B 6.80fF
C12641 sky130_fd_sc_hd__inv_1_53/Y sky130_fd_sc_hd__inv_1_53/A 0.08fF
C12642 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_17/a_1270_413# 0.00fF
C12643 sky130_fd_sc_hd__nor3_1_10/a_193_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12644 sky130_fd_sc_hd__nor3_1_6/a_193_297# DOUT[3] 0.00fF
C12645 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__inv_1_46/Y 0.00fF
C12646 sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C12647 sky130_fd_sc_hd__dfrtn_1_39/a_1217_47# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C12648 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# VDD 0.01fF
C12649 sky130_fd_sc_hd__nor3_1_5/A DOUT[9] 0.01fF
C12650 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# sky130_fd_sc_hd__inv_1_1/A 0.04fF
C12651 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C12652 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C12653 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__or3b_2_0/B 0.00fF
C12654 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__dfrtp_1_2/a_27_47# 0.00fF
C12655 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_2/a_193_47# 0.00fF
C12656 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_2/a_761_289# 0.00fF
C12657 sky130_fd_sc_hd__nor3_1_16/a_193_297# DOUT[16] 0.00fF
C12658 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__or2b_1_0/a_301_297# 0.00fF
C12659 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# sky130_fd_sc_hd__inv_1_47/A 0.01fF
C12660 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C12661 sky130_fd_sc_hd__nand3b_1_0/a_316_47# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C12662 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.01fF
C12663 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C12664 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.02fF
C12665 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C12666 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# RESET_COUNTERn 0.01fF
C12667 sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# sky130_fd_sc_hd__inv_1_38/A 0.00fF
C12668 DOUT[4] sky130_fd_sc_hd__dfrtn_1_35/a_805_47# 0.00fF
C12669 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# DOUT[21] 0.00fF
C12670 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_31/a_448_47# 0.00fF
C12671 VDD sky130_fd_sc_hd__inv_1_42/A 0.24fF
C12672 sky130_fd_sc_hd__nor3_1_4/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12673 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__or3b_2_0/a_176_21# 0.00fF
C12674 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__nor3_1_3/a_193_297# 0.00fF
C12675 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__nor3_1_3/a_109_297# 0.00fF
C12676 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C12677 sky130_fd_sc_hd__dfrtn_1_9/a_761_289# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C12678 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.03fF
C12679 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12680 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12681 sky130_fd_sc_hd__nand3b_1_1/a_316_47# VDD 0.00fF
C12682 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C12683 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# DOUT[11] 0.03fF
C12684 sky130_fd_sc_hd__dfrtn_1_4/a_761_289# VDD 0.05fF
C12685 sky130_fd_sc_hd__or3_1_0/a_183_297# VDD 0.00fF
C12686 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C12687 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# 0.00fF
C12688 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# 0.00fF
C12689 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__dfrtn_1_26/a_651_413# 0.00fF
C12690 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__dfrtn_1_28/a_193_47# 0.00fF
C12691 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# DOUT[3] 0.01fF
C12692 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C12693 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C12694 sky130_fd_sc_hd__dfrtn_1_32/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12695 sky130_fd_sc_hd__dfrtn_1_25/a_639_47# SEL_CONV_TIME[1] 0.00fF
C12696 sky130_fd_sc_hd__inv_1_1/Y RESET_COUNTERn 0.02fF
C12697 sky130_fd_sc_hd__nor3_2_1/a_281_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12698 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C12699 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_8/a_1270_413# 0.00fF
C12700 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# 0.00fF
C12701 sky130_fd_sc_hd__dfrtn_1_19/a_1108_47# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C12702 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C12703 sky130_fd_sc_hd__dfrtn_1_16/a_193_47# sky130_fd_sc_hd__dfrtn_1_16/a_1283_21# -0.00fF
C12704 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# sky130_fd_sc_hd__dfrtn_1_16/a_1108_47# -0.00fF
C12705 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12706 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# sky130_fd_sc_hd__inv_1_2/A 0.01fF
C12707 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# DOUT[3] 0.01fF
C12708 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__dfrtn_1_23/a_805_47# 0.00fF
C12709 sky130_fd_sc_hd__dfrtn_1_22/a_805_47# sky130_fd_sc_hd__dfrtn_1_23/a_27_47# 0.00fF
C12710 sky130_fd_sc_hd__dfrtn_1_31/a_1462_47# DONE 0.00fF
C12711 sky130_fd_sc_hd__dfrtn_1_21/a_543_47# sky130_fd_sc_hd__inv_1_30/Y 0.01fF
C12712 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C12713 sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C12714 sky130_fd_sc_hd__o311a_1_0/a_81_21# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C12715 sky130_fd_sc_hd__dfrtn_1_38/a_639_47# sky130_fd_sc_hd__inv_1_27/Y 0.00fF
C12716 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# sky130_fd_sc_hd__o311a_1_0/A3 0.01fF
C12717 sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# sky130_fd_sc_hd__dfrtn_1_21/a_193_47# -0.00fF
C12718 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C12719 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__inv_1_34/Y 0.01fF
C12720 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C12721 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_0/a_193_47# 0.59fF
C12722 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__dfrtn_1_16/a_1283_21# 0.00fF
C12723 sky130_fd_sc_hd__nor3_2_2/a_281_297# sky130_fd_sc_hd__dfrtn_1_16/a_543_47# 0.00fF
C12724 sky130_fd_sc_hd__mux4_2_0/a_193_369# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C12725 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__dfrtn_1_28/a_761_289# -0.00fF
C12726 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C12727 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__dfrtn_1_33/a_1217_47# 0.00fF
C12728 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__dfrtn_1_33/a_448_47# 0.00fF
C12729 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# VDD 0.17fF
C12730 sky130_fd_sc_hd__dfrtp_1_3/a_1270_413# RESET_COUNTERn 0.00fF
C12731 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_49/A 0.06fF
C12732 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_31/a_27_47# 0.00fF
C12733 sky130_fd_sc_hd__or3_1_0/X sky130_fd_sc_hd__or3_1_0/C 0.02fF
C12734 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__dfrtn_1_6/a_543_47# -0.00fF
C12735 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.00fF
C12736 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C12737 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.01fF
C12738 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.00fF
C12739 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C12740 sky130_fd_sc_hd__dfrtn_1_39/a_193_47# VDD 0.16fF
C12741 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12742 sky130_fd_sc_hd__dfrtn_1_25/a_1270_413# VDD 0.00fF
C12743 sky130_fd_sc_hd__dfrtn_1_25/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12744 sky130_fd_sc_hd__or2b_1_0/X sky130_fd_sc_hd__or3_1_0/X 0.00fF
C12745 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C12746 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__dfrtn_1_3/a_193_47# 0.00fF
C12747 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__dfrtn_1_3/a_543_47# 0.00fF
C12748 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_651_413# 0.00fF
C12749 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__dfrtn_1_3/a_27_47# 0.00fF
C12750 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__dfrtn_1_3/a_761_289# 0.00fF
C12751 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_3/a_448_47# 0.00fF
C12752 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C12753 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__nor3_1_5/a_109_297# 0.00fF
C12754 sky130_fd_sc_hd__dfrtn_1_18/a_193_47# VDD 0.12fF
C12755 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__inv_1_46/Y 0.00fF
C12756 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__dfrtn_1_25/a_27_47# 0.00fF
C12757 sky130_fd_sc_hd__dfrtn_1_20/a_651_413# sky130_fd_sc_hd__inv_1_35/Y 0.00fF
C12758 sky130_fd_sc_hd__inv_1_30/Y sky130_fd_sc_hd__inv_1_35/Y 0.01fF
C12759 sky130_fd_sc_hd__inv_1_11/A sky130_fd_sc_hd__inv_1_8/A 0.00fF
C12760 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__inv_1_5/Y 0.02fF
C12761 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# DOUT[2] 0.00fF
C12762 sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# 0.00fF
C12763 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# 0.00fF
C12764 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# 0.00fF
C12765 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C12766 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C12767 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C12768 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__inv_1_53/Y -0.02fF
C12769 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C12770 sky130_fd_sc_hd__dfrtn_1_24/a_448_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C12771 sky130_fd_sc_hd__dfrtn_1_42/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12772 sky130_fd_sc_hd__o211a_1_1/a_510_47# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C12773 sky130_fd_sc_hd__dfrtn_1_42/a_639_47# VDD -0.00fF
C12774 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# DOUT[14] 0.02fF
C12775 sky130_fd_sc_hd__o311a_1_0/a_266_47# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C12776 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C12777 sky130_fd_sc_hd__dfrtn_1_29/a_639_47# RESET_COUNTERn 0.00fF
C12778 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__nor3_1_4/a_109_297# 0.00fF
C12779 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_543_47# 0.00fF
C12780 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_761_289# 0.00fF
C12781 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C12782 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__inv_1_4/Y 0.04fF
C12783 sky130_fd_sc_hd__inv_1_13/Y sky130_fd_sc_hd__inv_1_5/A 0.00fF
C12784 sky130_fd_sc_hd__dfrtn_1_10/a_1270_413# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C12785 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C12786 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C12787 SEL_CONV_TIME[0] DOUT[21] 0.04fF
C12788 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_36/a_639_47# 0.00fF
C12789 sky130_fd_sc_hd__inv_1_32/A sky130_fd_sc_hd__inv_1_31/Y 0.23fF
C12790 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C12791 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C12792 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# sky130_fd_sc_hd__dfrtn_1_38/a_761_289# 0.00fF
C12793 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# sky130_fd_sc_hd__dfrtn_1_38/a_543_47# 0.00fF
C12794 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C12795 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__o311a_1_0/a_266_47# 0.00fF
C12796 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# DOUT[23] 0.00fF
C12797 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# VDD -0.00fF
C12798 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12799 sky130_fd_sc_hd__dfrtn_1_34/a_448_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C12800 sky130_fd_sc_hd__nor3_1_3/a_193_297# DOUT[7] 0.00fF
C12801 sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12802 sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# DOUT[11] 0.00fF
C12803 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_1/a_761_289# 0.00fF
C12804 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_1/a_543_47# 0.00fF
C12805 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_1/a_27_47# 0.00fF
C12806 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_1/a_193_47# 0.00fF
C12807 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# 0.00fF
C12808 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_639_47# 0.00fF
C12809 sky130_fd_sc_hd__o311a_1_0/a_266_297# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C12810 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.01fF
C12811 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# 0.00fF
C12812 sky130_fd_sc_hd__dfrtn_1_7/a_1217_47# DOUT[3] 0.00fF
C12813 sky130_fd_sc_hd__nor3_1_11/a_193_297# DOUT[19] 0.00fF
C12814 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C12815 sky130_fd_sc_hd__nor3_1_14/a_193_297# VDD 0.00fF
C12816 sky130_fd_sc_hd__mux4_2_0/a_288_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C12817 SLC_0/a_1235_416# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12818 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# SEL_CONV_TIME[1] 0.01fF
C12819 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# sky130_fd_sc_hd__dfrtn_1_7/a_761_289# -0.00fF
C12820 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_543_47# -0.00fF
C12821 sky130_fd_sc_hd__nor3_1_4/A VIN 0.00fF
C12822 sky130_fd_sc_hd__dfrtp_1_3/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12823 sky130_fd_sc_hd__dfrtn_1_16/a_1108_47# DOUT[15] 0.02fF
C12824 sky130_fd_sc_hd__nor3_1_18/a_109_297# sky130_fd_sc_hd__inv_1_39/Y 0.00fF
C12825 sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# sky130_fd_sc_hd__inv_1_43/A 0.03fF
C12826 sky130_fd_sc_hd__inv_1_28/A sky130_fd_sc_hd__or2_2_0/B 0.00fF
C12827 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__inv_1_28/Y 0.02fF
C12828 sky130_fd_sc_hd__dfrtn_1_7/a_1217_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C12829 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_5/Y 0.01fF
C12830 sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# DOUT[21] 0.01fF
C12831 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# RESET_COUNTERn 0.05fF
C12832 sky130_fd_sc_hd__dfrtn_1_26/a_761_289# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C12833 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__dfrtn_1_26/a_543_47# 0.00fF
C12834 sky130_fd_sc_hd__dfrtn_1_41/a_651_413# sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C12835 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# 0.00fF
C12836 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_639_47# 0.00fF
C12837 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# sky130_fd_sc_hd__dfrtn_1_7/a_651_413# 0.00fF
C12838 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# sky130_fd_sc_hd__dfrtn_1_7/a_193_47# 0.00fF
C12839 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# sky130_fd_sc_hd__dfrtn_1_7/a_761_289# 0.00fF
C12840 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# sky130_fd_sc_hd__dfrtn_1_7/a_27_47# 0.00fF
C12841 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C12842 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C12843 SEL_CONV_TIME[0] sky130_fd_sc_hd__o311a_1_0/A3 0.05fF
C12844 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_3/a_1217_47# 0.00fF
C12845 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__inv_1_11/A 0.07fF
C12846 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_0/a_1462_47# 0.00fF
C12847 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# DOUT[20] 0.01fF
C12848 sky130_fd_sc_hd__dfrtp_1_0/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12849 sky130_fd_sc_hd__nand3b_1_0/a_316_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C12850 sky130_fd_sc_hd__dfrtp_1_0/a_1217_47# VDD 0.00fF
C12851 sky130_fd_sc_hd__dfrtn_1_21/a_1270_413# RESET_COUNTERn 0.00fF
C12852 sky130_fd_sc_hd__nor3_2_3/C DOUT[0] 0.03fF
C12853 sky130_fd_sc_hd__nor3_1_1/a_193_297# DOUT[5] 0.00fF
C12854 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# RESET_COUNTERn 0.02fF
C12855 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# DOUT[20] 0.00fF
C12856 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# DOUT[7] 0.01fF
C12857 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# DOUT[6] 0.00fF
C12858 sky130_fd_sc_hd__inv_1_22/Y en 0.00fF
C12859 VDD sky130_fd_sc_hd__inv_1_2/Y 0.18fF
C12860 sky130_fd_sc_hd__dfrtn_1_22/a_805_47# RESET_COUNTERn 0.00fF
C12861 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C12862 sky130_fd_sc_hd__dfrtn_1_39/a_1462_47# VDD 0.00fF
C12863 CLK_REF sky130_fd_sc_hd__dfrtn_1_20/a_651_413# 0.00fF
C12864 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# 0.01fF
C12865 DOUT[9] DOUT[14] 0.00fF
C12866 sky130_fd_sc_hd__o2111a_2_0/a_386_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C12867 CLK_REF sky130_fd_sc_hd__inv_1_30/Y 0.03fF
C12868 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C12869 sky130_fd_sc_hd__inv_1_15/A VIN 0.12fF
C12870 sky130_fd_sc_hd__nor3_1_15/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12871 sky130_fd_sc_hd__dfrtn_1_30/a_651_413# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C12872 sky130_fd_sc_hd__nor3_1_16/a_109_297# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C12873 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# VDD 0.09fF
C12874 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_10/a_651_413# -0.00fF
C12875 sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# outb 0.00fF
C12876 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12877 sky130_fd_sc_hd__dfrtn_1_18/a_1462_47# VDD 0.00fF
C12878 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C12879 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C12880 DOUT[1] sky130_fd_sc_hd__nor3_2_3/A 0.01fF
C12881 sky130_fd_sc_hd__dfrtn_1_0/a_1462_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C12882 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# DOUT[14] 0.01fF
C12883 sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C12884 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C12885 sky130_fd_sc_hd__dfrtn_1_17/a_1270_413# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C12886 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# sky130_fd_sc_hd__inv_1_43/A 0.03fF
C12887 sky130_fd_sc_hd__dfrtn_1_16/a_1270_413# RESET_COUNTERn 0.00fF
C12888 sky130_fd_sc_hd__nor3_2_1/a_281_297# DOUT[0] 0.00fF
C12889 sky130_fd_sc_hd__dfrtn_1_8/a_1283_21# RESET_COUNTERn 0.01fF
C12890 sky130_fd_sc_hd__dfrtn_1_8/a_639_47# DOUT[21] 0.00fF
C12891 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# DOUT[14] 0.00fF
C12892 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__o211a_1_0/X 0.01fF
C12893 sky130_fd_sc_hd__dfrtn_1_9/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12894 VDD sky130_fd_sc_hd__dfrtn_1_9/a_639_47# 0.00fF
C12895 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# SEL_CONV_TIME[1] 0.02fF
C12896 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_20/a_639_47# -0.00fF
C12897 sky130_fd_sc_hd__dfrtn_1_20/a_761_289# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C12898 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C12899 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C12900 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# 0.00fF
C12901 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# 0.00fF
C12902 sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C12903 sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C12904 sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C12905 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# 0.00fF
C12906 sky130_fd_sc_hd__dfrtn_1_41/a_651_413# sky130_fd_sc_hd__dfrtn_1_38/a_639_47# 0.00fF
C12907 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__dfrtn_1_38/a_1462_47# 0.00fF
C12908 sky130_fd_sc_hd__dfrtn_1_32/a_543_47# sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C12909 sky130_fd_sc_hd__inv_1_39/Y sky130_fd_sc_hd__inv_1_40/A 0.00fF
C12910 sky130_fd_sc_hd__nor3_1_0/a_193_297# DOUT[18] 0.00fF
C12911 sky130_fd_sc_hd__dfrtn_1_19/a_1270_413# VDD 0.00fF
C12912 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_13/a_761_289# 0.00fF
C12913 sky130_fd_sc_hd__dfrtp_1_3/a_1217_47# DOUT[23] 0.00fF
C12914 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__or3_1_0/C 0.32fF
C12915 sky130_fd_sc_hd__dfrtn_1_26/a_761_289# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C12916 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C12917 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_18/a_1270_413# 0.00fF
C12918 sky130_fd_sc_hd__dfrtn_1_31/a_448_47# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C12919 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# 0.00fF
C12920 DOUT[4] sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# 0.00fF
C12921 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C12922 sky130_fd_sc_hd__nor3_1_2/a_193_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12923 sky130_fd_sc_hd__dfrtn_1_34/a_543_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C12924 sky130_fd_sc_hd__dfrtn_1_23/a_1217_47# RESET_COUNTERn 0.00fF
C12925 sky130_fd_sc_hd__dfrtn_1_22/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12926 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_9/Y 0.00fF
C12927 sky130_fd_sc_hd__dfrtn_1_7/a_805_47# DOUT[6] 0.00fF
C12928 sky130_fd_sc_hd__dfrtn_1_7/a_651_413# RESET_COUNTERn 0.00fF
C12929 sky130_fd_sc_hd__dfrtn_1_7/a_639_47# DOUT[7] 0.00fF
C12930 sky130_fd_sc_hd__dfrtn_1_7/a_1217_47# DOUT[20] 0.00fF
C12931 sky130_fd_sc_hd__dfrtn_1_10/a_1217_47# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C12932 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# VDD 0.21fF
C12933 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C12934 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_15/A 0.27fF
C12935 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C12936 sky130_fd_sc_hd__nor3_2_0/A sky130_fd_sc_hd__inv_1_8/A 0.11fF
C12937 sky130_fd_sc_hd__dfrtn_1_4/a_761_289# DOUT[3] 0.00fF
C12938 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C12939 sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.00fF
C12940 sky130_fd_sc_hd__inv_1_34/A VDD 0.34fF
C12941 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# DOUT[23] 0.00fF
C12942 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_0/a_805_47# -0.00fF
C12943 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# sky130_fd_sc_hd__dfrtn_1_0/a_639_47# -0.00fF
C12944 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C12945 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__dfrtn_1_35/a_761_289# -0.00fF
C12946 sky130_fd_sc_hd__dfrtp_1_1/a_448_47# CLK_REF 0.01fF
C12947 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C12948 sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C12949 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# DOUT[17] 0.00fF
C12950 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_1478_413# -0.00fF
C12951 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_0/a_750_97# -0.00fF
C12952 VDD sky130_fd_sc_hd__inv_1_39/Y 0.49fF
C12953 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C12954 sky130_fd_sc_hd__dfrtn_1_27/a_639_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C12955 sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# sky130_fd_sc_hd__dfrtn_1_27/a_543_47# 0.00fF
C12956 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# sky130_fd_sc_hd__dfrtn_1_27/a_651_413# 0.00fF
C12957 sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# sky130_fd_sc_hd__dfrtn_1_27/a_448_47# 0.00fF
C12958 sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C12959 sky130_fd_sc_hd__dfrtn_1_24/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12960 sky130_fd_sc_hd__dfrtn_1_24/a_1462_47# VDD 0.00fF
C12961 sky130_fd_sc_hd__dfrtn_1_16/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12962 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C12963 sky130_fd_sc_hd__dfrtn_1_8/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12964 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C12965 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# VDD 0.00fF
C12966 sky130_fd_sc_hd__dfrtn_1_36/a_761_289# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C12967 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__o211a_1_1/X 0.00fF
C12968 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C12969 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_31/a_651_413# 0.00fF
C12970 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C12971 sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# DOUT[14] 0.00fF
C12972 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_15/A 0.22fF
C12973 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_12/a_543_47# 0.01fF
C12974 DOUT[4] sky130_fd_sc_hd__dfrtn_1_32/a_193_47# 0.01fF
C12975 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C12976 sky130_fd_sc_hd__dfrtn_1_33/a_651_413# SEL_CONV_TIME[1] 0.00fF
C12977 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_543_47# 0.01fF
C12978 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C12979 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_17/a_761_289# 0.00fF
C12980 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C12981 sky130_fd_sc_hd__nor3_1_8/a_109_297# DOUT[14] 0.00fF
C12982 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# 0.00fF
C12983 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__dfrtn_1_14/a_193_47# 0.00fF
C12984 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_14/a_543_47# 0.00fF
C12985 sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# SEL_CONV_TIME[1] 0.00fF
C12986 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__dfrtn_1_42/a_193_47# 0.00fF
C12987 sky130_fd_sc_hd__nor3_2_2/a_281_297# sky130_fd_sc_hd__dfrtn_1_42/a_27_47# 0.00fF
C12988 sky130_fd_sc_hd__dfrtn_1_23/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C12989 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__inv_1_6/A 0.01fF
C12990 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__nor3_1_15/a_109_297# 0.00fF
C12991 sky130_fd_sc_hd__nor3_1_13/a_109_297# VDD 0.00fF
C12992 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C12993 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C12994 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# VDD 0.04fF
C12995 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C12996 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# sky130_fd_sc_hd__o221ai_1_0/a_493_297# 0.00fF
C12997 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C12998 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C12999 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# 0.00fF
C13000 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.00fF
C13001 sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13002 sky130_fd_sc_hd__dfrtn_1_11/a_805_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C13003 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C13004 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__nor3_1_3/a_109_297# 0.00fF
C13005 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13006 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# VDD 0.00fF
C13007 sky130_fd_sc_hd__nor3_1_7/a_109_297# VIN 0.00fF
C13008 sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# sky130_fd_sc_hd__dfrtn_1_23/a_193_47# 0.00fF
C13009 sky130_fd_sc_hd__dfrtn_1_42/a_1108_47# sky130_fd_sc_hd__dfrtn_1_23/a_27_47# 0.00fF
C13010 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C13011 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C13012 sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# SEL_CONV_TIME[1] 0.00fF
C13013 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C13014 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# RESET_COUNTERn 0.02fF
C13015 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13016 sky130_fd_sc_hd__nor3_2_3/B DOUT[7] 0.05fF
C13017 sky130_fd_sc_hd__dfrtn_1_11/a_1270_413# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C13018 sky130_fd_sc_hd__nor3_1_10/a_109_297# DOUT[8] 0.00fF
C13019 sky130_fd_sc_hd__nor3_1_10/a_193_297# DOUT[7] 0.00fF
C13020 sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C13021 sky130_fd_sc_hd__dfrtn_1_33/a_448_47# VDD 0.00fF
C13022 sky130_fd_sc_hd__dfrtn_1_3/a_761_289# RESET_COUNTERn 0.01fF
C13023 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# DOUT[3] 0.00fF
C13024 sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# VDD 0.00fF
C13025 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C13026 DOUT[23] DOUT[15] 0.72fF
C13027 sky130_fd_sc_hd__nor3_2_3/C DOUT[2] 0.17fF
C13028 sky130_fd_sc_hd__dfrtn_1_20/a_448_47# sky130_fd_sc_hd__inv_1_35/A 0.01fF
C13029 sky130_fd_sc_hd__nor3_1_0/a_193_297# DOUT[22] 0.00fF
C13030 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__nor3_1_4/a_193_297# 0.00fF
C13031 DOUT[4] sky130_fd_sc_hd__dfrtn_1_31/a_651_413# 0.00fF
C13032 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C13033 sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C13034 sky130_fd_sc_hd__dfrtn_1_30/a_639_47# sky130_fd_sc_hd__dfrtn_1_31/a_193_47# 0.00fF
C13035 sky130_fd_sc_hd__dfrtn_1_30/a_805_47# sky130_fd_sc_hd__dfrtn_1_31/a_27_47# 0.00fF
C13036 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_805_47# 0.00fF
C13037 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__dfrtn_1_31/a_639_47# 0.00fF
C13038 sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# sky130_fd_sc_hd__dfrtn_1_28/a_193_47# 0.00fF
C13039 sky130_fd_sc_hd__dfrtn_1_11/a_761_289# sky130_fd_sc_hd__inv_1_11/A 0.01fF
C13040 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# DOUT[14] 0.00fF
C13041 sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C13042 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C13043 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__dfrtn_1_17/a_1270_413# 0.00fF
C13044 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__or2_2_0/B 0.15fF
C13045 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# HEADER_0/a_508_138# 0.00fF
C13046 DOUT[13] sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C13047 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__inv_1_33/A 0.00fF
C13048 sky130_fd_sc_hd__inv_1_46/Y VDD 0.17fF
C13049 sky130_fd_sc_hd__o211a_1_1/a_215_47# sky130_fd_sc_hd__dfrtn_1_17/a_651_413# 0.00fF
C13050 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__dfrtn_1_17/a_639_47# 0.00fF
C13051 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# DOUT[17] 0.01fF
C13052 sky130_fd_sc_hd__dfrtn_1_34/a_1270_413# SEL_CONV_TIME[1] 0.00fF
C13053 sky130_fd_sc_hd__nor3_1_14/a_193_297# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C13054 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_448_47# 0.00fF
C13055 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C13056 sky130_fd_sc_hd__dfrtn_1_24/a_448_47# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C13057 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# 0.00fF
C13058 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# sky130_fd_sc_hd__dfrtn_1_29/a_543_47# 0.00fF
C13059 sky130_fd_sc_hd__dfrtn_1_25/a_805_47# SEL_CONV_TIME[0] 0.00fF
C13060 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C13061 sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# VDD 0.10fF
C13062 sky130_fd_sc_hd__inv_1_22/Y VIN 0.13fF
C13063 sky130_fd_sc_hd__dfrtn_1_33/a_761_289# sky130_fd_sc_hd__inv_1_45/A 0.01fF
C13064 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# 0.00fF
C13065 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__inv_1_12/A 0.03fF
C13066 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# sky130_fd_sc_hd__dfrtn_1_11/a_543_47# 0.00fF
C13067 sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# 0.00fF
C13068 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_11/a_639_47# 0.00fF
C13069 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# 0.00fF
C13070 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__dfrtn_1_11/a_651_413# 0.00fF
C13071 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_805_47# 0.00fF
C13072 SEL_CONV_TIME[3] RESET_COUNTERn 0.01fF
C13073 sky130_fd_sc_hd__nor3_2_3/a_27_297# VDD 0.07fF
C13074 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C13075 sky130_fd_sc_hd__inv_1_7/Y RESET_COUNTERn 0.04fF
C13076 sky130_fd_sc_hd__dfrtn_1_42/a_761_289# DOUT[15] 0.00fF
C13077 DOUT[4] sky130_fd_sc_hd__dfrtn_1_32/a_1462_47# 0.00fF
C13078 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/a_448_47# -0.00fF
C13079 sky130_fd_sc_hd__dfrtn_1_7/a_448_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C13080 sky130_fd_sc_hd__inv_1_2/Y DOUT[3] 0.47fF
C13081 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# 0.00fF
C13082 sky130_fd_sc_hd__dfrtn_1_12/a_805_47# sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# 0.00fF
C13083 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# 0.00fF
C13084 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__dfrtn_1_34/a_27_47# 0.00fF
C13085 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# -0.00fF
C13086 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_37/a_448_47# -0.00fF
C13087 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_14/a_639_47# 0.00fF
C13088 sky130_fd_sc_hd__dfrtn_1_28/a_651_413# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C13089 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C13090 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13091 sky130_fd_sc_hd__dfrtn_1_26/a_448_47# VDD 0.01fF
C13092 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__inv_1_47/Y 0.00fF
C13093 sky130_fd_sc_hd__nor3_1_0/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13094 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C13095 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_2/Y 0.06fF
C13096 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# DOUT[14] 0.00fF
C13097 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__o2111a_2_0/a_386_47# 0.00fF
C13098 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__o2111a_2_0/a_80_21# 0.00fF
C13099 sky130_fd_sc_hd__inv_1_6/A DOUT[8] 0.10fF
C13100 sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13101 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C13102 sky130_fd_sc_hd__dfrtn_1_34/a_651_413# VDD 0.01fF
C13103 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C13104 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13105 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# 0.00fF
C13106 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__dfrtn_1_30/a_651_413# 0.00fF
C13107 sky130_fd_sc_hd__or2b_1_0/a_301_297# sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# 0.00fF
C13108 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_8/a_193_47# 0.01fF
C13109 sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C13110 sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C13111 sky130_fd_sc_hd__dfrtn_1_23/a_448_47# sky130_fd_sc_hd__inv_1_40/Y 0.02fF
C13112 sky130_fd_sc_hd__dfrtn_1_28/a_651_413# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C13113 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# -0.00fF
C13114 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_3/a_543_47# -0.00fF
C13115 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__inv_1_17/A 0.00fF
C13116 sky130_fd_sc_hd__o221ai_1_0/a_295_297# SEL_CONV_TIME[0] 0.00fF
C13117 sky130_fd_sc_hd__o2111a_2_0/a_566_47# SEL_CONV_TIME[1] 0.01fF
C13118 SEL_CONV_TIME[2] RESET_COUNTERn 0.18fF
C13119 sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# RESET_COUNTERn 0.02fF
C13120 sky130_fd_sc_hd__dfrtn_1_25/a_639_47# DOUT[21] 0.00fF
C13121 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_6/a_805_47# 0.00fF
C13122 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__or2_2_0/X 0.26fF
C13123 sky130_fd_sc_hd__nand3b_1_1/Y sky130_fd_sc_hd__inv_1_33/A 0.01fF
C13124 sky130_fd_sc_hd__inv_1_4/A DOUT[6] 0.00fF
C13125 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__inv_1_32/Y 0.01fF
C13126 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C13127 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C13128 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C13129 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__o211a_1_1/a_297_297# 0.00fF
C13130 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.00fF
C13131 sky130_fd_sc_hd__dfrtp_1_0/a_1283_21# DOUT[15] 0.00fF
C13132 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C13133 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C13134 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_26/a_761_289# 0.01fF
C13135 sky130_fd_sc_hd__inv_1_40/Y DOUT[21] 0.00fF
C13136 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__or2b_1_0/X 0.01fF
C13137 DOUT[4] sky130_fd_sc_hd__dfrtn_1_29/a_761_289# 0.00fF
C13138 DOUT[13] sky130_fd_sc_hd__or3b_2_0/a_388_297# 0.00fF
C13139 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__inv_1_43/A 0.02fF
C13140 sky130_fd_sc_hd__dfrtn_1_7/a_651_413# HEADER_0/a_508_138# 0.00fF
C13141 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C13142 sky130_fd_sc_hd__dfrtn_1_28/a_193_47# SEL_CONV_TIME[1] 0.00fF
C13143 sky130_fd_sc_hd__dfrtn_1_40/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13144 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# VDD 0.00fF
C13145 sky130_fd_sc_hd__mux4_2_0/a_600_345# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C13146 sky130_fd_sc_hd__dfrtn_1_42/a_1108_47# RESET_COUNTERn 0.02fF
C13147 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# SEL_CONV_TIME[3] 0.00fF
C13148 sky130_fd_sc_hd__inv_1_36/A sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C13149 sky130_fd_sc_hd__nor3_1_12/a_193_297# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C13150 sky130_fd_sc_hd__dfrtn_1_0/a_1462_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C13151 sky130_fd_sc_hd__dfrtn_1_34/a_639_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C13152 sky130_fd_sc_hd__nor3_1_16/a_193_297# RESET_COUNTERn 0.00fF
C13153 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C13154 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# 0.00fF
C13155 sky130_fd_sc_hd__dfrtn_1_0/a_639_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C13156 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__or3_1_0/C 0.01fF
C13157 sky130_fd_sc_hd__mux4_2_0/a_193_369# sky130_fd_sc_hd__mux4_2_0/a_288_47# -0.00fF
C13158 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtp_1_3/a_761_289# 0.00fF
C13159 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtp_1_3/a_651_413# 0.00fF
C13160 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtp_1_3/a_543_47# 0.00fF
C13161 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_448_47# 0.00fF
C13162 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C13163 sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C13164 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13165 sky130_fd_sc_hd__o2111a_2_0/a_458_47# VDD 0.00fF
C13166 DOUT[13] sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# 0.00fF
C13167 sky130_fd_sc_hd__nor3_1_20/a_109_297# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C13168 HEADER_0/a_508_138# RESET_COUNTERn 0.03fF
C13169 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# DOUT[20] 0.00fF
C13170 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# RESET_COUNTERn 0.00fF
C13171 sky130_fd_sc_hd__dfrtn_1_17/a_639_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C13172 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C13173 sky130_fd_sc_hd__dfrtn_1_4/a_639_47# RESET_COUNTERn 0.00fF
C13174 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# SEL_CONV_TIME[0] 0.00fF
C13175 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__dfrtn_1_34/a_543_47# 0.00fF
C13176 sky130_fd_sc_hd__or2b_1_0/a_301_297# sky130_fd_sc_hd__dfrtn_1_34/a_193_47# 0.00fF
C13177 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C13178 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__nor3_1_3/a_109_297# 0.00fF
C13179 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__nor3_1_3/a_193_297# 0.00fF
C13180 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13181 SLC_0/a_264_22# RESET_COUNTERn 0.03fF
C13182 sky130_fd_sc_hd__dfrtn_1_31/a_1283_21# sky130_fd_sc_hd__inv_1_49/A 0.03fF
C13183 DOUT[13] sky130_fd_sc_hd__dfrtn_1_31/a_761_289# 0.00fF
C13184 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_27_47# 0.00fF
C13185 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# SEL_CONV_TIME[2] 0.01fF
C13186 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_29/a_761_289# 0.00fF
C13187 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__or3b_2_0/B 0.00fF
C13188 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# VDD 0.17fF
C13189 sky130_fd_sc_hd__inv_1_26/A lc_out 0.02fF
C13190 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_193_47# -0.00fF
C13191 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__o2111a_2_0/X 0.01fF
C13192 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C13193 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__nor3_1_13/a_109_297# 0.00fF
C13194 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C13195 sky130_fd_sc_hd__dfrtn_1_14/a_651_413# VDD 0.00fF
C13196 sky130_fd_sc_hd__dfrtn_1_12/a_1462_47# sky130_fd_sc_hd__dfrtn_1_0/a_27_47# 0.00fF
C13197 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_0/a_1462_47# 0.00fF
C13198 sky130_fd_sc_hd__dfrtn_1_7/a_543_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C13199 sky130_fd_sc_hd__inv_1_23/A DOUT[10] 0.00fF
C13200 sky130_fd_sc_hd__dfrtn_1_37/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13201 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# DOUT[3] 0.00fF
C13202 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C13203 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# RESET_COUNTERn 0.00fF
C13204 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__inv_1_8/Y 0.01fF
C13205 DOUT[10] RESET_COUNTERn 0.00fF
C13206 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# -0.00fF
C13207 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C13208 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# 0.00fF
C13209 sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13210 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_8/a_1462_47# 0.00fF
C13211 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C13212 sky130_fd_sc_hd__inv_1_2/Y DOUT[20] 0.01fF
C13213 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C13214 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C13215 sky130_fd_sc_hd__dfrtn_1_39/a_1270_413# RESET_COUNTERn 0.00fF
C13216 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C13217 sky130_fd_sc_hd__dfrtn_1_22/a_448_47# sky130_fd_sc_hd__inv_1_39/Y 0.01fF
C13218 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__inv_1_13/A 0.01fF
C13219 sky130_fd_sc_hd__dfrtn_1_42/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C13220 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# DOUT[21] 0.01fF
C13221 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__inv_1_42/A 0.01fF
C13222 sky130_fd_sc_hd__dfrtp_1_3/a_1217_47# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C13223 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__nor3_1_3/a_193_297# 0.00fF
C13224 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__nand2_1_1/a_113_47# 0.00fF
C13225 sky130_fd_sc_hd__dfrtn_1_18/a_1270_413# RESET_COUNTERn -0.00fF
C13226 VDD sky130_fd_sc_hd__mux4_1_0/X 0.31fF
C13227 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__dfrtn_1_25/a_761_289# 0.00fF
C13228 sky130_fd_sc_hd__or3_1_0/a_111_297# sky130_fd_sc_hd__dfrtn_1_25/a_193_47# 0.00fF
C13229 sky130_fd_sc_hd__or3_1_0/a_183_297# sky130_fd_sc_hd__dfrtn_1_25/a_27_47# 0.00fF
C13230 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# 0.00fF
C13231 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__nor3_2_2/A 0.01fF
C13232 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C13233 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__inv_1_13/A 0.40fF
C13234 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__inv_1_36/A 0.01fF
C13235 sky130_fd_sc_hd__dfrtn_1_4/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13236 SEL_CONV_TIME[2] SEL_CONV_TIME[3] 0.05fF
C13237 sky130_fd_sc_hd__dfrtn_1_30/a_761_289# SEL_CONV_TIME[0] 0.02fF
C13238 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# 0.00fF
C13239 sky130_fd_sc_hd__dfrtn_1_3/a_651_413# sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C13240 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C13241 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__dfrtn_1_7/a_27_47# 0.00fF
C13242 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__dfrtn_1_7/a_193_47# 0.00fF
C13243 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C13244 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# DOUT[3] 0.00fF
C13245 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# VDD 0.05fF
C13246 DOUT[11] sky130_fd_sc_hd__nor3_2_3/C 0.23fF
C13247 sky130_fd_sc_hd__inv_1_26/A sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C13248 sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# RESET_COUNTERn 0.02fF
C13249 sky130_fd_sc_hd__nor3_2_0/A sky130_fd_sc_hd__inv_1_15/A 0.00fF
C13250 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_193_47# 0.00fF
C13251 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_27_47# 0.00fF
C13252 sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# sky130_fd_sc_hd__dfrtp_1_3/a_651_413# 0.00fF
C13253 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C13254 sky130_fd_sc_hd__dfrtn_1_19/a_1283_21# RESET_COUNTERn 0.00fF
C13255 CLK_REF sky130_fd_sc_hd__dfrtn_1_17/a_1270_413# 0.00fF
C13256 sky130_fd_sc_hd__inv_1_15/A DOUT[17] 0.01fF
C13257 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C13258 sky130_fd_sc_hd__o311a_1_0/a_266_297# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C13259 sky130_fd_sc_hd__mux4_2_0/a_600_345# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C13260 sky130_fd_sc_hd__nor3_1_17/a_109_297# RESET_COUNTERn 0.00fF
C13261 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C13262 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# -0.29fF
C13263 sky130_fd_sc_hd__dfrtp_1_0/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13264 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_543_47# 0.00fF
C13265 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C13266 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_4/a_761_289# 0.00fF
C13267 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C13268 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__inv_1_43/Y 0.04fF
C13269 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__inv_1_8/A 0.01fF
C13270 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_448_47# -0.00fF
C13271 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_651_413# -0.00fF
C13272 sky130_fd_sc_hd__dfrtn_1_21/a_1270_413# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C13273 sky130_fd_sc_hd__or3b_2_0/a_472_297# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C13274 sky130_fd_sc_hd__dfrtn_1_35/a_543_47# sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# 0.00fF
C13275 sky130_fd_sc_hd__dfrtn_1_35/a_448_47# sky130_fd_sc_hd__dfrtn_1_36/a_761_289# 0.00fF
C13276 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_1270_413# 0.00fF
C13277 sky130_fd_sc_hd__dfrtn_1_35/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_651_413# 0.00fF
C13278 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# 0.00fF
C13279 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# 0.00fF
C13280 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_1217_47# 0.00fF
C13281 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C13282 sky130_fd_sc_hd__dfrtn_1_28/a_1217_47# VDD 0.00fF
C13283 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C13284 sky130_fd_sc_hd__nand3b_1_1/Y sky130_fd_sc_hd__o2111a_2_0/X 0.10fF
C13285 sky130_fd_sc_hd__dfrtn_1_27/a_193_47# sky130_fd_sc_hd__inv_1_43/A 0.03fF
C13286 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C13287 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_37/a_448_47# 0.01fF
C13288 sky130_fd_sc_hd__dfrtn_1_0/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C13289 sky130_fd_sc_hd__dfrtn_1_9/a_651_413# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C13290 sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# VDD 0.08fF
C13291 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# VDD 0.22fF
C13292 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__inv_1_15/A 0.24fF
C13293 sky130_fd_sc_hd__nor3_1_13/a_109_297# sky130_fd_sc_hd__dfrtn_1_8/a_27_47# 0.00fF
C13294 sky130_fd_sc_hd__inv_1_14/A sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C13295 sky130_fd_sc_hd__or3_1_0/X RESET_COUNTERn 0.00fF
C13296 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__nand3b_1_1/Y 0.01fF
C13297 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C13298 sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# sky130_fd_sc_hd__inv_1_14/A 0.03fF
C13299 sky130_fd_sc_hd__mux4_1_0/a_668_97# SEL_CONV_TIME[1] 0.00fF
C13300 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# 0.00fF
C13301 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C13302 sky130_fd_sc_hd__nand3b_1_0/a_232_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C13303 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_38/a_1270_413# 0.00fF
C13304 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C13305 DOUT[9] sky130_fd_sc_hd__dfrtn_1_3/a_651_413# 0.00fF
C13306 sky130_fd_sc_hd__nor3_1_3/a_193_297# VIN 0.00fF
C13307 sky130_fd_sc_hd__nor3_1_5/a_109_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13308 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C13309 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_14/a_543_47# 0.01fF
C13310 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C13311 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C13312 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_24/a_27_47# 0.00fF
C13313 sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# sky130_fd_sc_hd__inv_1_32/Y 0.00fF
C13314 sky130_fd_sc_hd__dfrtn_1_20/a_639_47# VDD 0.00fF
C13315 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_193_47# -0.33fF
C13316 sky130_fd_sc_hd__dfrtn_1_25/a_1217_47# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C13317 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# sky130_fd_sc_hd__or2_2_0/A 0.01fF
C13318 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# RESET_COUNTERn 0.04fF
C13319 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__inv_1_32/Y 0.03fF
C13320 sky130_fd_sc_hd__dfrtn_1_9/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13321 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# SEL_CONV_TIME[1] 0.00fF
C13322 sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# sky130_fd_sc_hd__inv_1_32/Y 0.01fF
C13323 CLK_REF sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.37fF
C13324 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_2/a_543_47# 0.00fF
C13325 DOUT[1] sky130_fd_sc_hd__dfrtn_1_36/a_639_47# 0.00fF
C13326 DOUT[4] sky130_fd_sc_hd__dfrtn_1_8/a_1270_413# 0.00fF
C13327 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__inv_1_31/A 0.00fF
C13328 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_4/a_448_47# 0.00fF
C13329 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_12/a_543_47# -0.00fF
C13330 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_12/a_761_289# -0.00fF
C13331 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_26/a_805_47# 0.00fF
C13332 DOUT[9] sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C13333 sky130_fd_sc_hd__dfrtn_1_16/a_448_47# DOUT[2] 0.00fF
C13334 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# sky130_fd_sc_hd__dfrtn_1_42/a_805_47# -0.00fF
C13335 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# 0.00fF
C13336 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_543_47# 0.00fF
C13337 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__dfrtn_1_13/a_193_47# 0.00fF
C13338 sky130_fd_sc_hd__o221ai_1_0/a_213_123# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13339 sky130_fd_sc_hd__nor3_1_18/a_109_297# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C13340 DOUT[9] sky130_fd_sc_hd__dfrtn_1_4/a_543_47# 0.00fF
C13341 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# DOUT[11] 0.00fF
C13342 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__dfrtp_1_0/a_761_289# -0.00fF
C13343 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C13344 sky130_fd_sc_hd__mux4_1_0/a_193_47# VDD 0.00fF
C13345 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C13346 sky130_fd_sc_hd__dfrtn_1_10/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13347 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C13348 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C13349 sky130_fd_sc_hd__o211a_1_0/a_297_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13350 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_19/a_651_413# 0.00fF
C13351 sky130_fd_sc_hd__o211a_1_0/a_510_47# VDD -0.00fF
C13352 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# 0.00fF
C13353 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# VIN 0.04fF
C13354 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__inv_1_51/Y 0.01fF
C13355 sky130_fd_sc_hd__dfrtp_1_0/a_805_47# DOUT[23] 0.00fF
C13356 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# 0.01fF
C13357 sky130_fd_sc_hd__or2_2_0/a_39_297# sky130_fd_sc_hd__or2_2_0/A 0.01fF
C13358 sky130_fd_sc_hd__dfrtn_1_27/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_651_413# -0.00fF
C13359 sky130_fd_sc_hd__nor3_1_13/a_193_297# DOUT[21] 0.00fF
C13360 sky130_fd_sc_hd__nor3_2_2/A RESET_COUNTERn 0.32fF
C13361 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C13362 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_11/a_651_413# 0.00fF
C13363 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C13364 sky130_fd_sc_hd__mux4_2_0/a_1064_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C13365 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_4/a_805_47# 0.00fF
C13366 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# DOUT[7] 0.00fF
C13367 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# DOUT[20] 0.00fF
C13368 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# 0.00fF
C13369 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__dfrtn_1_4/a_651_413# 0.00fF
C13370 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# sky130_fd_sc_hd__dfrtn_1_4/a_543_47# 0.00fF
C13371 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# sky130_fd_sc_hd__dfrtn_1_4/a_448_47# 0.00fF
C13372 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# RESET_COUNTERn 0.03fF
C13373 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# -0.00fF
C13374 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__dfrtn_1_29/a_448_47# 0.00fF
C13375 sky130_fd_sc_hd__dfrtn_1_39/a_1270_413# SEL_CONV_TIME[2] 0.00fF
C13376 sky130_fd_sc_hd__inv_1_33/A sky130_fd_sc_hd__inv_1_32/Y 0.13fF
C13377 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C13378 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C13379 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_39/a_27_47# 0.01fF
C13380 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__o311a_1_0/a_266_47# 0.00fF
C13381 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__o311a_1_0/a_585_47# 0.00fF
C13382 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__inv_1_45/A 0.18fF
C13383 sky130_fd_sc_hd__inv_1_53/A RESET_COUNTERn 0.15fF
C13384 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# 0.00fF
C13385 sky130_fd_sc_hd__dfrtn_1_39/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C13386 DOUT[1] sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# 0.00fF
C13387 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__dfrtn_1_14/a_27_47# 0.00fF
C13388 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C13389 sky130_fd_sc_hd__dfrtn_1_33/a_761_289# RESET_COUNTERn 0.01fF
C13390 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# DOUT[19] 0.00fF
C13391 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C13392 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__mux4_2_0/a_600_345# 0.00fF
C13393 sky130_fd_sc_hd__dfrtn_1_27/a_1462_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C13394 sky130_fd_sc_hd__nor3_1_1/a_193_297# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C13395 sky130_fd_sc_hd__dfrtn_1_24/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13396 sky130_fd_sc_hd__dfrtn_1_35/a_1217_47# VDD 0.00fF
C13397 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13398 sky130_fd_sc_hd__nor3_2_1/a_27_297# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C13399 sky130_fd_sc_hd__dfrtn_1_12/a_1217_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C13400 sky130_fd_sc_hd__dfrtn_1_30/a_651_413# RESET_COUNTERn 0.00fF
C13401 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.01fF
C13402 sky130_fd_sc_hd__nor3_2_1/a_27_297# sky130_fd_sc_hd__o211a_1_0/a_215_47# 0.00fF
C13403 SLC_0/a_1235_416# sky130_fd_sc_hd__inv_1_26/A 0.00fF
C13404 sky130_fd_sc_hd__nor3_1_11/a_109_297# VDD 0.00fF
C13405 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C13406 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.00fF
C13407 sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# SEL_CONV_TIME[0] 0.00fF
C13408 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C13409 sky130_fd_sc_hd__dfrtn_1_18/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# -0.00fF
C13410 sky130_fd_sc_hd__dfrtn_1_18/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# -0.00fF
C13411 sky130_fd_sc_hd__dfrtn_1_18/a_761_289# sky130_fd_sc_hd__dfrtn_1_18/a_543_47# -0.00fF
C13412 sky130_fd_sc_hd__mux4_2_0/a_872_316# SEL_CONV_TIME[1] 0.00fF
C13413 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# DOUT[19] 0.00fF
C13414 sky130_fd_sc_hd__dfrtn_1_27/a_805_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C13415 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C13416 sky130_fd_sc_hd__dfrtn_1_34/a_639_47# SEL_CONV_TIME[0] 0.00fF
C13417 sky130_fd_sc_hd__dfrtp_1_1/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C13418 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__inv_1_31/Y 0.20fF
C13419 sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# VDD 0.00fF
C13420 sky130_fd_sc_hd__dfrtn_1_23/a_1462_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C13421 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_30/a_639_47# 0.00fF
C13422 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C13423 sky130_fd_sc_hd__inv_1_37/A sky130_fd_sc_hd__inv_1_40/A 0.00fF
C13424 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C13425 sky130_fd_sc_hd__dfrtn_1_16/a_543_47# sky130_fd_sc_hd__inv_1_25/A 0.00fF
C13426 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# SLC_0/a_264_22# 0.00fF
C13427 sky130_fd_sc_hd__dfrtp_1_0/a_1108_47# SLC_0/a_1235_416# 0.00fF
C13428 sky130_fd_sc_hd__or3_1_0/X SEL_CONV_TIME[3] 0.06fF
C13429 SLC_0/a_438_293# out 0.01fF
C13430 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# RESET_COUNTERn 0.31fF
C13431 sky130_fd_sc_hd__dfrtn_1_14/a_761_289# DOUT[18] 0.00fF
C13432 sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# SEL_CONV_TIME[1] 0.00fF
C13433 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C13434 CLK_REF sky130_fd_sc_hd__dfrtp_1_3/a_1217_47# 0.00fF
C13435 sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C13436 sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# sky130_fd_sc_hd__or2_2_0/a_121_297# 0.00fF
C13437 sky130_fd_sc_hd__nor3_2_1/a_27_297# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C13438 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# 0.00fF
C13439 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# 0.00fF
C13440 sky130_fd_sc_hd__dfrtn_1_7/a_651_413# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C13441 sky130_fd_sc_hd__dfrtn_1_8/a_1270_413# outb 0.00fF
C13442 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_10/a_543_47# 0.02fF
C13443 DOUT[9] sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# 0.00fF
C13444 sky130_fd_sc_hd__dfrtn_1_10/a_805_47# sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# 0.00fF
C13445 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# 0.00fF
C13446 sky130_fd_sc_hd__o311a_1_0/a_266_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13447 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__inv_1_33/A 0.04fF
C13448 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_1_24/A 0.01fF
C13449 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_12/a_1270_413# 0.00fF
C13450 sky130_fd_sc_hd__dfrtn_1_7/a_639_47# VIN 0.00fF
C13451 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C13452 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C13453 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C13454 sky130_fd_sc_hd__mux4_2_0/a_193_47# VDD 0.00fF
C13455 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# out 0.00fF
C13456 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C13457 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__inv_1_44/A 0.01fF
C13458 sky130_fd_sc_hd__inv_1_4/Y RESET_COUNTERn 0.03fF
C13459 sky130_fd_sc_hd__dfrtn_1_18/a_27_47# sky130_fd_sc_hd__inv_1_33/A 0.02fF
C13460 sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# SEL_CONV_TIME[1] 0.00fF
C13461 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_2/a_761_289# 0.01fF
C13462 sky130_fd_sc_hd__inv_1_42/Y RESET_COUNTERn 0.02fF
C13463 sky130_fd_sc_hd__dfrtn_1_26/a_761_289# RESET_COUNTERn 0.02fF
C13464 sky130_fd_sc_hd__dfrtn_1_34/a_1217_47# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C13465 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C13466 sky130_fd_sc_hd__dfrtp_1_1/a_448_47# sky130_fd_sc_hd__nor3_2_1/a_281_297# 0.00fF
C13467 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__nor3_2_1/a_27_297# 0.00fF
C13468 sky130_fd_sc_hd__or3_1_0/X SEL_CONV_TIME[2] 0.00fF
C13469 sky130_fd_sc_hd__or3b_2_0/X sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13470 sky130_fd_sc_hd__dfrtn_1_33/a_543_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C13471 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C13472 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.01fF
C13473 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C13474 sky130_fd_sc_hd__dfrtn_1_35/a_448_47# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C13475 sky130_fd_sc_hd__dfrtn_1_16/a_193_47# sky130_fd_sc_hd__nor3_2_3/A 0.54fF
C13476 sky130_fd_sc_hd__dfrtn_1_34/a_543_47# RESET_COUNTERn 0.00fF
C13477 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13478 sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# VDD 0.07fF
C13479 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13480 sky130_fd_sc_hd__dfrtp_1_2/a_805_47# RESET_COUNTERn 0.00fF
C13481 sky130_fd_sc_hd__dfrtn_1_35/a_1108_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C13482 sky130_fd_sc_hd__nor3_1_20/a_193_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13483 sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13484 sky130_fd_sc_hd__dfrtn_1_41/a_805_47# VDD 0.00fF
C13485 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C13486 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# DOUT[2] 0.00fF
C13487 VDD sky130_fd_sc_hd__inv_1_37/A 1.80fF
C13488 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C13489 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# 0.00fF
C13490 sky130_fd_sc_hd__dfrtn_1_8/a_543_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C13491 sky130_fd_sc_hd__dfrtn_1_21/a_193_47# sky130_fd_sc_hd__dfrtn_1_19/a_1270_413# 0.00fF
C13492 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_35/a_27_47# 0.01fF
C13493 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_39/a_1217_47# 0.00fF
C13494 sky130_fd_sc_hd__o211a_1_1/X sky130_fd_sc_hd__dfrtp_1_1/D 0.01fF
C13495 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# DONE 0.00fF
C13496 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__mux4_1_0/a_277_47# 0.11fF
C13497 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_30/a_805_47# 0.00fF
C13498 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C13499 sky130_fd_sc_hd__dfrtn_1_28/a_761_289# SEL_CONV_TIME[0] 0.00fF
C13500 sky130_fd_sc_hd__mux4_2_0/a_1060_369# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C13501 sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13502 sky130_fd_sc_hd__dfrtn_1_27/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C13503 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C13504 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C13505 sky130_fd_sc_hd__dfrtn_1_27/a_543_47# VDD 0.04fF
C13506 sky130_fd_sc_hd__dfrtn_1_34/a_1270_413# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C13507 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_18/a_543_47# 0.02fF
C13508 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__dfrtn_1_1/a_193_47# 0.00fF
C13509 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__dfrtn_1_1/a_761_289# 0.00fF
C13510 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# RESET_COUNTERn 0.01fF
C13511 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C13512 sky130_fd_sc_hd__inv_1_3/Y sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C13513 sky130_fd_sc_hd__o211a_1_1/a_215_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C13514 sky130_fd_sc_hd__dfrtn_1_36/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_761_289# -0.00fF
C13515 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_543_47# -0.00fF
C13516 sky130_fd_sc_hd__inv_1_53/A SEL_CONV_TIME[3] 0.13fF
C13517 sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C13518 sky130_fd_sc_hd__dfrtn_1_29/a_639_47# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C13519 sky130_fd_sc_hd__o2111a_2_0/a_566_47# DOUT[21] 0.00fF
C13520 sky130_fd_sc_hd__nor3_1_3/a_109_297# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C13521 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C13522 sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# RESET_COUNTERn 0.00fF
C13523 sky130_fd_sc_hd__dfrtn_1_26/a_543_47# sky130_fd_sc_hd__inv_1_43/Y 0.01fF
C13524 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_21/a_193_47# 0.29fF
C13525 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C13526 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# VDD 0.06fF
C13527 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13528 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_639_47# 0.00fF
C13529 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C13530 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C13531 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_448_47# 0.00fF
C13532 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C13533 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C13534 sky130_fd_sc_hd__nor3_2_3/B VIN 0.07fF
C13535 sky130_fd_sc_hd__nor3_1_10/a_193_297# VIN 0.00fF
C13536 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# 0.00fF
C13537 sky130_fd_sc_hd__dfrtp_1_3/a_1108_47# sky130_fd_sc_hd__or2_2_0/B 0.01fF
C13538 sky130_fd_sc_hd__nor3_1_15/a_109_297# DOUT[1] 0.00fF
C13539 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13540 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C13541 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C13542 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# VDD 0.01fF
C13543 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# 0.00fF
C13544 sky130_fd_sc_hd__dfrtn_1_39/a_1217_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C13545 sky130_fd_sc_hd__dfrtn_1_17/a_651_413# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C13546 sky130_fd_sc_hd__nor3_1_5/A VDD 1.24fF
C13547 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_1/a_27_47# 0.01fF
C13548 sky130_fd_sc_hd__dfrtn_1_28/a_193_47# DOUT[21] 0.01fF
C13549 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13550 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__nor3_1_1/a_109_297# 0.00fF
C13551 sky130_fd_sc_hd__dfrtn_1_33/a_1108_47# DOUT[23] 0.00fF
C13552 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_805_47# -0.00fF
C13553 sky130_fd_sc_hd__inv_1_53/A SEL_CONV_TIME[2] 0.45fF
C13554 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_5/Y 0.09fF
C13555 sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# DOUT[5] 0.00fF
C13556 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# DOUT[14] 0.00fF
C13557 sky130_fd_sc_hd__dfrtn_1_14/a_543_47# RESET_COUNTERn 0.01fF
C13558 sky130_fd_sc_hd__mux4_1_0/a_193_413# SEL_CONV_TIME[0] 0.00fF
C13559 sky130_fd_sc_hd__dfrtn_1_28/a_1108_47# sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C13560 sky130_fd_sc_hd__dfrtn_1_18/a_1217_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C13561 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__inv_1_47/Y 0.00fF
C13562 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C13563 sky130_fd_sc_hd__dfrtn_1_42/a_1108_47# sky130_fd_sc_hd__nor3_2_2/A 0.02fF
C13564 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_34/a_448_47# 0.00fF
C13565 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__dfrtp_1_3/a_651_413# 0.00fF
C13566 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# sky130_fd_sc_hd__dfrtp_1_3/a_1270_413# 0.00fF
C13567 sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C13568 sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C13569 sky130_fd_sc_hd__dfrtn_1_16/a_1462_47# sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C13570 sky130_fd_sc_hd__dfrtn_1_33/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13571 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C13572 sky130_fd_sc_hd__dfrtn_1_36/a_448_47# sky130_fd_sc_hd__inv_1_40/A 0.00fF
C13573 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# VIN 0.00fF
C13574 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__nand3b_1_1/a_232_47# 0.00fF
C13575 sky130_fd_sc_hd__dfrtn_1_14/a_761_289# DOUT[22] 0.00fF
C13576 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# 0.01fF
C13577 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# 0.01fF
C13578 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_37/a_761_289# 0.00fF
C13579 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_37/a_448_47# 0.00fF
C13580 sky130_fd_sc_hd__dfrtn_1_40/a_1270_413# sky130_fd_sc_hd__dfrtn_1_37/a_193_47# 0.00fF
C13581 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_37/a_651_413# 0.00fF
C13582 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_37/a_639_47# 0.00fF
C13583 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__dfrtn_1_37/a_27_47# 0.00fF
C13584 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__dfrtn_1_34/a_27_47# 0.00fF
C13585 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__dfrtn_1_34/a_193_47# 0.00fF
C13586 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C13587 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13588 sky130_fd_sc_hd__inv_1_42/Y SEL_CONV_TIME[3] 0.08fF
C13589 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C13590 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# 0.00fF
C13591 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C13592 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__dfrtn_1_2/a_761_289# 0.00fF
C13593 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_639_47# 0.00fF
C13594 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C13595 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__dfrtn_1_2/a_651_413# 0.00fF
C13596 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_25/a_27_47# 0.00fF
C13597 sky130_fd_sc_hd__dfrtn_1_34/a_1462_47# DONE 0.00fF
C13598 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C13599 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C13600 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# -0.00fF
C13601 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# -0.00fF
C13602 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# 0.00fF
C13603 sky130_fd_sc_hd__dfrtn_1_42/a_543_47# DOUT[2] 0.00fF
C13604 sky130_fd_sc_hd__dfrtn_1_27/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13605 DOUT[9] sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# 0.00fF
C13606 sky130_fd_sc_hd__dfrtn_1_38/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13607 sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C13608 DOUT[1] sky130_fd_sc_hd__dfrtn_1_22/a_651_413# 0.00fF
C13609 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_34/a_27_47# 0.01fF
C13610 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__inv_1_31/Y 0.17fF
C13611 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_41/a_543_47# 0.01fF
C13612 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.01fF
C13613 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13614 sky130_fd_sc_hd__or3_1_0/C sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C13615 sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# DOUT[23] 0.00fF
C13616 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C13617 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# DOUT[19] 0.01fF
C13618 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# DOUT[14] 0.00fF
C13619 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# 0.01fF
C13620 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__dfrtn_1_15/a_27_47# 0.00fF
C13621 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_448_47# 0.00fF
C13622 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C13623 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_15/a_543_47# 0.00fF
C13624 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# 0.00fF
C13625 sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C13626 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C13627 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C13628 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C13629 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C13630 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C13631 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# 0.00fF
C13632 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C13633 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__inv_1_54/Y 0.00fF
C13634 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# sky130_fd_sc_hd__nor3_1_0/a_109_297# 0.00fF
C13635 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# sky130_fd_sc_hd__nor3_1_0/a_193_297# 0.00fF
C13636 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C13637 sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C13638 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C13639 sky130_fd_sc_hd__dfrtn_1_36/a_448_47# VDD 0.01fF
C13640 sky130_fd_sc_hd__dfrtn_1_12/a_761_289# sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# 0.00fF
C13641 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_651_413# 0.00fF
C13642 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__dfrtn_1_13/a_193_47# 0.00fF
C13643 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# 0.00fF
C13644 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C13645 sky130_fd_sc_hd__inv_1_9/A sky130_fd_sc_hd__nor3_2_3/C 1.09fF
C13646 sky130_fd_sc_hd__inv_1_26/A DOUT[2] 0.00fF
C13647 sky130_fd_sc_hd__dfrtn_1_0/a_805_47# DOUT[18] 0.00fF
C13648 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# 0.00fF
C13649 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__or2b_1_0/X 0.01fF
C13650 sky130_fd_sc_hd__nor3_2_3/a_281_297# sky130_fd_sc_hd__dfrtn_1_42/a_27_47# 0.00fF
C13651 sky130_fd_sc_hd__nor3_2_3/a_27_297# sky130_fd_sc_hd__dfrtn_1_42/a_193_47# 0.00fF
C13652 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# 0.00fF
C13653 sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13654 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_13/a_193_47# 0.00fF
C13655 sky130_fd_sc_hd__dfrtn_1_0/a_1270_413# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C13656 sky130_fd_sc_hd__nor3_1_13/a_109_297# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C13657 sky130_fd_sc_hd__nor3_1_11/a_109_297# DOUT[3] 0.00fF
C13658 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_27/a_805_47# 0.00fF
C13659 sky130_fd_sc_hd__dfrtn_1_34/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13660 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C13661 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13662 sky130_fd_sc_hd__dfrtn_1_28/a_1462_47# DOUT[21] 0.00fF
C13663 sky130_fd_sc_hd__dfrtn_1_28/a_651_413# RESET_COUNTERn 0.00fF
C13664 sky130_fd_sc_hd__dfrtn_1_30/a_1270_413# sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C13665 sky130_fd_sc_hd__nor3_1_11/a_109_297# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C13666 sky130_fd_sc_hd__nor3_1_3/a_109_297# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C13667 sky130_fd_sc_hd__mux4_1_0/a_834_97# SEL_CONV_TIME[0] 0.00fF
C13668 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# 0.00fF
C13669 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__nor3_2_3/B 0.13fF
C13670 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# RESET_COUNTERn 0.01fF
C13671 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13672 sky130_fd_sc_hd__dfrtn_1_35/a_193_47# DOUT[21] 0.01fF
C13673 HEADER_0/a_508_138# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C13674 sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C13675 sky130_fd_sc_hd__dfrtn_1_23/a_761_289# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C13676 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C13677 DOUT[4] sky130_fd_sc_hd__dfrtn_1_24/a_193_47# 0.00fF
C13678 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_543_47# 0.00fF
C13679 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_761_289# 0.00fF
C13680 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_39/a_27_47# 0.00fF
C13681 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_30/a_27_47# 0.02fF
C13682 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# SEL_CONV_TIME[2] 0.00fF
C13683 sky130_fd_sc_hd__inv_1_31/Y sky130_fd_sc_hd__inv_1_33/A 0.01fF
C13684 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# VIN 0.00fF
C13685 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__inv_1_43/A 0.01fF
C13686 sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# 0.00fF
C13687 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__dfrtn_1_21/a_761_289# -0.00fF
C13688 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C13689 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# 0.00fF
C13690 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C13691 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C13692 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C13693 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C13694 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_448_47# 0.00fF
C13695 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C13696 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C13697 sky130_fd_sc_hd__dfrtn_1_32/a_448_47# sky130_fd_sc_hd__inv_1_9/A 0.00fF
C13698 sky130_fd_sc_hd__inv_1_47/A RESET_COUNTERn 0.39fF
C13699 sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# RESET_COUNTERn 0.00fF
C13700 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# SEL_CONV_TIME[0] 0.00fF
C13701 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__inv_1_29/Y 0.00fF
C13702 DOUT[1] sky130_fd_sc_hd__dfrtn_1_23/a_1270_413# 0.00fF
C13703 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_543_47# 0.00fF
C13704 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C13705 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.00fF
C13706 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_761_289# 0.00fF
C13707 sky130_fd_sc_hd__dfrtn_1_18/a_448_47# DOUT[2] 0.00fF
C13708 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# sky130_fd_sc_hd__inv_1_25/A 0.02fF
C13709 sky130_fd_sc_hd__dfrtn_1_32/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C13710 sky130_fd_sc_hd__dfrtn_1_32/a_761_289# VDD 0.05fF
C13711 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_25/a_1217_47# 0.00fF
C13712 VDD sky130_fd_sc_hd__nor3_1_19/Y 0.87fF
C13713 DOUT[9] DOUT[19] 0.02fF
C13714 sky130_fd_sc_hd__dfrtn_1_22/a_1462_47# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C13715 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# DOUT[11] 0.01fF
C13716 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C13717 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_448_47# -0.00fF
C13718 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# -0.00fF
C13719 sky130_fd_sc_hd__dfrtn_1_36/a_193_47# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C13720 DOUT[16] sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C13721 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__nand3b_1_0/Y 0.00fF
C13722 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_38/a_543_47# 0.00fF
C13723 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# sky130_fd_sc_hd__inv_1_52/Y 0.55fF
C13724 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C13725 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_34/a_1217_47# 0.00fF
C13726 sky130_fd_sc_hd__dfrtn_1_31/a_639_47# SEL_CONV_TIME[1] 0.00fF
C13727 sky130_fd_sc_hd__mux4_1_0/a_750_97# RESET_COUNTERn 0.01fF
C13728 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.01fF
C13729 sky130_fd_sc_hd__dfrtn_1_10/a_805_47# RESET_COUNTERn 0.00fF
C13730 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C13731 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_28/a_27_47# 0.01fF
C13732 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_24/a_193_47# 0.00fF
C13733 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_448_47# 0.00fF
C13734 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_31/a_651_413# 0.00fF
C13735 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_19/a_1217_47# 0.00fF
C13736 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# DOUT[19] 0.00fF
C13737 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C13738 sky130_fd_sc_hd__inv_1_41/Y sky130_fd_sc_hd__inv_1_48/A 0.01fF
C13739 sky130_fd_sc_hd__nor3_1_14/a_193_297# outb 0.00fF
C13740 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# 0.00fF
C13741 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# 0.00fF
C13742 sky130_fd_sc_hd__dfrtn_1_17/a_805_47# VDD 0.00fF
C13743 sky130_fd_sc_hd__dfrtn_1_28/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C13744 sky130_fd_sc_hd__dfrtn_1_3/a_1462_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C13745 VDD DOUT[14] 2.17fF
C13746 sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13747 sky130_fd_sc_hd__dfrtn_1_0/a_761_289# sky130_fd_sc_hd__nor3_1_0/a_109_297# 0.00fF
C13748 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_37/A 0.01fF
C13749 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# sky130_fd_sc_hd__nor3_1_0/a_193_297# 0.00fF
C13750 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13751 sky130_fd_sc_hd__dfrtn_1_32/a_27_47# sky130_fd_sc_hd__dfrtn_1_32/a_448_47# -0.00fF
C13752 sky130_fd_sc_hd__dfrtn_1_32/a_193_47# sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# -0.00fF
C13753 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# 0.00fF
C13754 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__dfrtn_1_24/a_27_47# 0.00fF
C13755 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__nor3_1_5/A 0.05fF
C13756 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# 0.00fF
C13757 sky130_fd_sc_hd__dfrtn_1_22/a_448_47# sky130_fd_sc_hd__inv_1_37/A 0.01fF
C13758 sky130_fd_sc_hd__dfrtn_1_3/a_805_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C13759 DOUT[4] sky130_fd_sc_hd__dfrtn_1_30/a_27_47# 0.00fF
C13760 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__dfrtn_1_30/a_761_289# -0.00fF
C13761 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__dfrtn_1_30/a_543_47# -0.00fF
C13762 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C13763 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_448_47# 0.00fF
C13764 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C13765 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C13766 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C13767 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfrtn_1_41/a_543_47# 0.01fF
C13768 sky130_fd_sc_hd__nor3_1_10/a_109_297# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C13769 sky130_fd_sc_hd__dfrtn_1_31/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13770 sky130_fd_sc_hd__dfrtn_1_31/a_1270_413# VDD 0.00fF
C13771 sky130_fd_sc_hd__mux4_2_0/a_397_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C13772 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C13773 sky130_fd_sc_hd__dfrtn_1_38/a_543_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C13774 sky130_fd_sc_hd__dfrtn_1_28/a_543_47# sky130_fd_sc_hd__inv_1_42/A 0.01fF
C13775 sky130_fd_sc_hd__mux4_2_0/a_1060_369# SEL_CONV_TIME[0] 0.00fF
C13776 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__mux4_1_0/X 0.01fF
C13777 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__inv_1_15/A 0.01fF
C13778 sky130_fd_sc_hd__dfrtn_1_35/a_651_413# RESET_COUNTERn 0.00fF
C13779 sky130_fd_sc_hd__dfrtn_1_0/a_1217_47# RESET_COUNTERn 0.00fF
C13780 sky130_fd_sc_hd__inv_1_11/A sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C13781 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# sky130_fd_sc_hd__dfrtn_1_31/a_448_47# -0.00fF
C13782 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_651_413# -0.00fF
C13783 sky130_fd_sc_hd__dfrtn_1_29/a_805_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C13784 sky130_fd_sc_hd__nor3_1_11/a_109_297# DOUT[20] 0.00fF
C13785 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# DOUT[3] 0.00fF
C13786 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# 0.00fF
C13787 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# 0.00fF
C13788 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_39/a_1462_47# 0.00fF
C13789 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_39/a_1217_47# 0.00fF
C13790 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_14/a_27_47# 0.00fF
C13791 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# RESET_COUNTERn 0.04fF
C13792 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_761_289# 0.00fF
C13793 sky130_fd_sc_hd__dfrtp_1_3/a_543_47# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C13794 sky130_fd_sc_hd__dfrtp_1_3/a_761_289# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C13795 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_543_47# 0.00fF
C13796 sky130_fd_sc_hd__dfrtn_1_4/a_448_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C13797 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_19/a_639_47# 0.00fF
C13798 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_19/a_805_47# 0.00fF
C13799 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__inv_1_31/A 0.00fF
C13800 sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# sky130_fd_sc_hd__inv_1_35/Y 0.00fF
C13801 sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# SEL_CONV_TIME[0] 0.00fF
C13802 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C13803 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_38/a_805_47# 0.00fF
C13804 sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C13805 sky130_fd_sc_hd__dfrtn_1_34/a_651_413# sky130_fd_sc_hd__o221ai_1_0/a_493_297# 0.00fF
C13806 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C13807 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_18/a_1462_47# 0.00fF
C13808 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_18/a_1217_47# 0.00fF
C13809 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_18/a_1270_413# 0.00fF
C13810 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C13811 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_18/a_651_413# 0.00fF
C13812 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# 0.00fF
C13813 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_40/a_193_47# 0.00fF
C13814 sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13815 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C13816 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__dfrtn_1_29/a_543_47# 0.00fF
C13817 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C13818 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__dfrtn_1_29/a_761_289# 0.00fF
C13819 sky130_fd_sc_hd__inv_1_48/A sky130_fd_sc_hd__inv_1_49/A 0.01fF
C13820 sky130_fd_sc_hd__dfrtn_1_32/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13821 sky130_fd_sc_hd__dfrtn_1_10/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13822 sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C13823 DOUT[13] sky130_fd_sc_hd__inv_1_50/Y 0.22fF
C13824 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C13825 sky130_fd_sc_hd__dfrtp_1_3/a_761_289# VDD 0.04fF
C13826 sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C13827 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_1/a_448_47# -0.00fF
C13828 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# -0.00fF
C13829 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# SEL_CONV_TIME[1] 0.01fF
C13830 sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C13831 sky130_fd_sc_hd__nor3_1_5/A DOUT[5] 0.00fF
C13832 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_21/a_805_47# 0.00fF
C13833 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__or3_1_0/X 0.01fF
C13834 sky130_fd_sc_hd__o311a_1_0/a_266_297# RESET_COUNTERn 0.00fF
C13835 sky130_fd_sc_hd__dfrtp_1_3/a_639_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C13836 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C13837 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C13838 sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# SEL_CONV_TIME[0] 0.00fF
C13839 sky130_fd_sc_hd__mux4_2_0/a_872_316# DOUT[21] 0.00fF
C13840 sky130_fd_sc_hd__mux4_2_0/a_288_47# RESET_COUNTERn 0.00fF
C13841 sky130_fd_sc_hd__or2_2_0/a_39_297# RESET_COUNTERn 0.02fF
C13842 sky130_fd_sc_hd__dfrtn_1_23/a_651_413# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C13843 sky130_fd_sc_hd__dfrtn_1_25/a_1217_47# sky130_fd_sc_hd__dfrtn_1_28/a_27_47# 0.00fF
C13844 sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# sky130_fd_sc_hd__dfrtn_1_28/a_448_47# 0.00fF
C13845 sky130_fd_sc_hd__nor3_1_18/a_193_297# sky130_fd_sc_hd__nor3_2_2/a_27_297# 0.00fF
C13846 sky130_fd_sc_hd__nor3_1_18/a_109_297# sky130_fd_sc_hd__nor3_2_2/a_281_297# 0.00fF
C13847 CLK_REF sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C13848 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_36/a_448_47# 0.00fF
C13849 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C13850 sky130_fd_sc_hd__nor3_1_15/a_109_297# sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# 0.00fF
C13851 sky130_fd_sc_hd__nor3_1_15/a_193_297# sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.00fF
C13852 sky130_fd_sc_hd__nor3_1_4/A DOUT[8] 0.00fF
C13853 sky130_fd_sc_hd__nor3_1_8/a_109_297# DOUT[19] 0.00fF
C13854 sky130_fd_sc_hd__nor3_1_15/a_193_297# sky130_fd_sc_hd__inv_1_9/A 0.00fF
C13855 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C13856 sky130_fd_sc_hd__dfrtn_1_42/a_639_47# sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C13857 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_6/A 0.02fF
C13858 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# RESET_COUNTERn 0.14fF
C13859 sky130_fd_sc_hd__dfrtn_1_4/a_651_413# DOUT[11] 0.00fF
C13860 sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13861 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# -0.00fF
C13862 sky130_fd_sc_hd__dfrtn_1_35/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13863 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# VDD 0.00fF
C13864 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C13865 sky130_fd_sc_hd__dfrtn_1_41/a_448_47# RESET_COUNTERn 0.00fF
C13866 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_34/a_651_413# 0.00fF
C13867 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__or2_2_0/B 0.00fF
C13868 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__nor3_2_1/a_281_297# 0.00fF
C13869 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__nor3_2_1/a_27_297# 0.00fF
C13870 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C13871 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# VDD 0.05fF
C13872 DOUT[4] sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# 0.00fF
C13873 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C13874 sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# sky130_fd_sc_hd__inv_1_8/A 0.01fF
C13875 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C13876 sky130_fd_sc_hd__dfrtn_1_19/a_1270_413# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C13877 sky130_fd_sc_hd__dfrtn_1_3/a_651_413# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C13878 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__o211a_1_1/a_215_47# 0.00fF
C13879 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.00fF
C13880 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__o211a_1_1/a_510_47# 0.00fF
C13881 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__o211a_1_1/a_297_297# 0.00fF
C13882 sky130_fd_sc_hd__dfrtn_1_20/a_761_289# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.00fF
C13883 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.00fF
C13884 sky130_fd_sc_hd__dfrtn_1_25/a_1217_47# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C13885 sky130_fd_sc_hd__dfrtn_1_32/a_651_413# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C13886 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__o211a_1_1/X 0.00fF
C13887 sky130_fd_sc_hd__dfrtn_1_23/a_761_289# sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C13888 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C13889 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_761_289# 0.00fF
C13890 sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# DOUT[21] 0.00fF
C13891 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__inv_1_53/A 0.02fF
C13892 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C13893 CLK_REF sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# 0.00fF
C13894 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_1/a_651_413# 0.00fF
C13895 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__inv_1_38/A 0.02fF
C13896 sky130_fd_sc_hd__inv_1_39/A sky130_fd_sc_hd__nor3_2_3/B 0.30fF
C13897 sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C13898 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# sky130_fd_sc_hd__inv_1_12/A 0.01fF
C13899 sky130_fd_sc_hd__nor3_2_1/A DOUT[23] 0.01fF
C13900 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__dfrtn_1_25/a_761_289# 0.00fF
C13901 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_25/a_651_413# 0.00fF
C13902 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__dfrtn_1_25/a_543_47# 0.00fF
C13903 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__nor3_1_2/a_193_297# 0.00fF
C13904 sky130_fd_sc_hd__dfrtp_1_3/a_639_47# sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# 0.00fF
C13905 sky130_fd_sc_hd__dfrtp_1_3/a_761_289# sky130_fd_sc_hd__dfrtn_1_17/a_1462_47# 0.00fF
C13906 sky130_fd_sc_hd__dfrtp_1_3/a_543_47# sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# 0.00fF
C13907 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_32/a_761_289# 0.00fF
C13908 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C13909 sky130_fd_sc_hd__nor3_1_15/a_193_297# sky130_fd_sc_hd__dfrtn_1_32/a_27_47# 0.00fF
C13910 sky130_fd_sc_hd__nor3_1_10/a_109_297# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C13911 sky130_fd_sc_hd__dfrtn_1_12/a_805_47# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C13912 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.01fF
C13913 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.00fF
C13914 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__mux4_2_0/a_600_345# 0.00fF
C13915 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# sky130_fd_sc_hd__mux4_2_0/a_193_369# 0.00fF
C13916 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C13917 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# sky130_fd_sc_hd__mux4_2_0/a_372_413# 0.00fF
C13918 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13919 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__inv_1_7/A 0.01fF
C13920 sky130_fd_sc_hd__dfrtn_1_4/a_543_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C13921 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13922 sky130_fd_sc_hd__inv_1_14/A DOUT[11] 0.02fF
C13923 sky130_fd_sc_hd__inv_1_18/Y sky130_fd_sc_hd__inv_1_22/Y 0.01fF
C13924 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C13925 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# 0.00fF
C13926 sky130_fd_sc_hd__dfrtn_1_4/a_805_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C13927 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C13928 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C13929 sky130_fd_sc_hd__o2111a_2_0/a_458_47# sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# 0.00fF
C13930 sky130_fd_sc_hd__o2111a_2_0/a_386_47# sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# 0.00fF
C13931 sky130_fd_sc_hd__a221oi_4_0/a_27_297# SEL_CONV_TIME[0] 0.01fF
C13932 sky130_fd_sc_hd__dfrtp_1_3/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13933 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# RESET_COUNTERn 0.02fF
C13934 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__inv_1_28/A 0.00fF
C13935 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C13936 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# 0.00fF
C13937 sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C13938 sky130_fd_sc_hd__dfrtn_1_22/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13939 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C13940 sky130_fd_sc_hd__dfrtn_1_22/a_1283_21# VDD 0.09fF
C13941 DOUT[1] sky130_fd_sc_hd__dfrtn_1_42/a_761_289# 0.00fF
C13942 sky130_fd_sc_hd__dfrtn_1_12/a_761_289# RESET_COUNTERn 0.01fF
C13943 sky130_fd_sc_hd__dfrtn_1_20/a_761_289# sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# 0.01fF
C13944 sky130_fd_sc_hd__dfrtn_1_20/a_639_47# sky130_fd_sc_hd__dfrtn_1_21/a_193_47# 0.00fF
C13945 sky130_fd_sc_hd__dfrtn_1_41/a_651_413# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C13946 sky130_fd_sc_hd__or2_2_0/B DOUT[23] 0.02fF
C13947 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C13948 sky130_fd_sc_hd__dfrtn_1_28/a_448_47# sky130_fd_sc_hd__inv_1_48/A 0.01fF
C13949 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# 0.00fF
C13950 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C13951 DOUT[4] sky130_fd_sc_hd__dfrtn_1_34/a_651_413# 0.00fF
C13952 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# DOUT[2] 0.01fF
C13953 sky130_fd_sc_hd__nor3_1_13/a_109_297# outb 0.00fF
C13954 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C13955 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__dfrtn_1_6/a_193_47# 0.00fF
C13956 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__dfrtn_1_6/a_27_47# 0.00fF
C13957 sky130_fd_sc_hd__nor3_1_2/a_193_297# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C13958 sky130_fd_sc_hd__dfrtp_1_1/a_639_47# sky130_fd_sc_hd__dfrtp_1_1/D 0.00fF
C13959 sky130_fd_sc_hd__nand3b_1_0/a_232_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C13960 sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# sky130_fd_sc_hd__inv_1_40/A 0.02fF
C13961 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__dfrtp_1_1/a_27_47# 0.00fF
C13962 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# -0.00fF
C13963 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C13964 sky130_fd_sc_hd__dfrtn_1_11/a_1462_47# RESET_COUNTERn 0.00fF
C13965 sky130_fd_sc_hd__dfrtn_1_8/a_761_289# sky130_fd_sc_hd__inv_1_9/A 0.01fF
C13966 sky130_fd_sc_hd__o311a_1_0/a_266_297# SEL_CONV_TIME[3] 0.00fF
C13967 sky130_fd_sc_hd__nor3_2_0/A sky130_fd_sc_hd__nor3_2_3/B 0.26fF
C13968 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_10/a_651_413# 0.00fF
C13969 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_761_289# 0.00fF
C13970 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C13971 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C13972 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# DOUT[23] 0.00fF
C13973 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# DOUT[19] 0.00fF
C13974 sky130_fd_sc_hd__dfrtn_1_8/a_651_413# DOUT[12] 0.00fF
C13975 sky130_fd_sc_hd__nor3_1_0/a_193_297# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C13976 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C13977 sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# sky130_fd_sc_hd__nor3_2_0/A 0.01fF
C13978 sky130_fd_sc_hd__mux4_2_0/a_288_47# SEL_CONV_TIME[3] 0.01fF
C13979 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__inv_1_12/A 0.01fF
C13980 sky130_fd_sc_hd__dfrtn_1_16/a_761_289# VDD 0.05fF
C13981 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.03fF
C13982 SLC_0/a_438_293# sky130_fd_sc_hd__o211a_1_0/a_79_21# 0.00fF
C13983 sky130_fd_sc_hd__o211a_1_0/a_297_297# sky130_fd_sc_hd__inv_1_26/A 0.00fF
C13984 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13985 sky130_fd_sc_hd__nor3_2_3/B DOUT[17] 0.04fF
C13986 sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C13987 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C13988 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_1108_47# -0.00fF
C13989 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__dfrtp_1_3/a_448_47# -0.00fF
C13990 sky130_fd_sc_hd__nand3b_1_1/Y sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C13991 sky130_fd_sc_hd__inv_1_14/A sky130_fd_sc_hd__nor3_1_5/a_109_297# 0.00fF
C13992 VDD SEL_CONV_TIME[0] 5.29fF
C13993 CLK_REF sky130_fd_sc_hd__dfrtn_1_19/a_651_413# 0.00fF
C13994 sky130_fd_sc_hd__nor3_2_2/a_281_297# VDD 0.04fF
C13995 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__inv_1_1/A 0.01fF
C13996 sky130_fd_sc_hd__dfrtn_1_20/a_1462_47# sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.00fF
C13997 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_20/a_27_47# 0.01fF
C13998 sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# sky130_fd_sc_hd__dfrtn_1_18/a_639_47# 0.00fF
C13999 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C14000 sky130_fd_sc_hd__inv_1_6/Y sky130_fd_sc_hd__inv_1_6/A 0.03fF
C14001 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__dfrtn_1_29/a_448_47# 0.00fF
C14002 sky130_fd_sc_hd__dfrtn_1_18/a_448_47# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C14003 sky130_fd_sc_hd__inv_1_12/A sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C14004 SEL_CONV_TIME[1] DOUT[21] 0.67fF
C14005 sky130_fd_sc_hd__dfrtp_1_0/a_1283_21# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C14006 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C14007 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_13/A 0.00fF
C14008 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_34/a_651_413# 0.00fF
C14009 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_40/a_193_47# -0.06fF
C14010 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# sky130_fd_sc_hd__o211a_1_0/a_510_47# 0.00fF
C14011 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# sky130_fd_sc_hd__o211a_1_0/a_79_21# 0.00fF
C14012 sky130_fd_sc_hd__dfrtn_1_23/a_1462_47# sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C14013 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# sky130_fd_sc_hd__dfrtn_1_36/a_639_47# 0.00fF
C14014 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C14015 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# -0.00fF
C14016 sky130_fd_sc_hd__dfrtn_1_27/a_805_47# RESET_COUNTERn 0.00fF
C14017 DOUT[3] DOUT[14] 0.00fF
C14018 sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C14019 sky130_fd_sc_hd__dfrtn_1_35/a_1217_47# sky130_fd_sc_hd__inv_1_38/A 0.00fF
C14020 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C14021 sky130_fd_sc_hd__mux4_2_0/a_288_47# SEL_CONV_TIME[2] 0.01fF
C14022 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__nor3_1_0/a_109_297# 0.00fF
C14023 sky130_fd_sc_hd__nor3_1_11/a_193_297# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C14024 sky130_fd_sc_hd__dfrtn_1_9/a_448_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C14025 sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# VDD 0.07fF
C14026 sky130_fd_sc_hd__dfrtn_1_23/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14027 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14028 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_35/a_1283_21# 0.00fF
C14029 sky130_fd_sc_hd__dfrtn_1_30/a_1270_413# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C14030 sky130_fd_sc_hd__nor3_2_0/a_281_297# sky130_fd_sc_hd__dfrtn_1_12/a_651_413# 0.00fF
C14031 sky130_fd_sc_hd__inv_1_2/A DOUT[14] 0.47fF
C14032 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__dfrtn_1_34/a_448_47# -0.00fF
C14033 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# -0.00fF
C14034 DOUT[13] sky130_fd_sc_hd__dfrtn_1_30/a_448_47# 0.01fF
C14035 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C14036 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C14037 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_38/a_543_47# 0.00fF
C14038 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C14039 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C14040 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_448_47# 0.00fF
C14041 sky130_fd_sc_hd__dfrtn_1_38/a_639_47# DOUT[2] 0.00fF
C14042 sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# sky130_fd_sc_hd__mux4_2_0/a_600_345# 0.00fF
C14043 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# sky130_fd_sc_hd__mux4_2_0/a_1281_47# 0.00fF
C14044 sky130_fd_sc_hd__dfrtn_1_37/a_1462_47# sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C14045 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# sky130_fd_sc_hd__mux4_2_0/a_1064_47# 0.00fF
C14046 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# VDD 0.07fF
C14047 sky130_fd_sc_hd__mux4_2_0/a_1064_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14048 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# sky130_fd_sc_hd__inv_1_32/A 0.01fF
C14049 sky130_fd_sc_hd__dfrtn_1_36/a_761_289# RESET_COUNTERn 0.03fF
C14050 sky130_fd_sc_hd__dfrtn_1_36/a_651_413# DOUT[21] 0.00fF
C14051 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__inv_1_5/Y 0.01fF
C14052 DOUT[4] sky130_fd_sc_hd__dfrtn_1_28/a_27_47# 0.00fF
C14053 sky130_fd_sc_hd__dfrtp_1_0/a_1283_21# sky130_fd_sc_hd__or2_2_0/B 0.01fF
C14054 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# RESET_COUNTERn 0.00fF
C14055 SEL_CONV_TIME[1] sky130_fd_sc_hd__o311a_1_0/A3 0.02fF
C14056 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C14057 sky130_fd_sc_hd__inv_1_28/Y sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14058 sky130_fd_sc_hd__dfrtn_1_9/a_639_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C14059 sky130_fd_sc_hd__dfrtn_1_14/a_651_413# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C14060 sky130_fd_sc_hd__dfrtn_1_33/a_543_47# sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# 0.00fF
C14061 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C14062 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C14063 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# VDD 0.01fF
C14064 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# 0.00fF
C14065 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# -0.00fF
C14066 sky130_fd_sc_hd__nor3_1_12/a_109_297# sky130_fd_sc_hd__dfrtn_1_8/a_651_413# 0.00fF
C14067 sky130_fd_sc_hd__nor3_1_12/a_193_297# sky130_fd_sc_hd__dfrtn_1_8/a_448_47# 0.00fF
C14068 sky130_fd_sc_hd__dfrtn_1_11/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14069 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C14070 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C14071 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__dfrtn_1_25/a_651_413# 0.00fF
C14072 sky130_fd_sc_hd__dfrtn_1_21/a_805_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C14073 sky130_fd_sc_hd__dfrtn_1_18/a_639_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C14074 sky130_fd_sc_hd__o2111a_2_0/a_386_47# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C14075 sky130_fd_sc_hd__nor3_1_7/a_193_297# DOUT[7] 0.00fF
C14076 sky130_fd_sc_hd__dfrtn_1_27/a_761_289# DOUT[23] 0.00fF
C14077 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# 0.00fF
C14078 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# 0.00fF
C14079 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# 0.00fF
C14080 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/a_805_47# 0.00fF
C14081 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__mux4_2_0/a_1064_47# 0.00fF
C14082 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# DOUT[0] 0.00fF
C14083 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.00fF
C14084 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_761_289# 0.00fF
C14085 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C14086 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_543_47# 0.01fF
C14087 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.00fF
C14088 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__nor3_1_4/a_193_297# 0.00fF
C14089 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C14090 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__dfrtn_1_13/a_761_289# 0.00fF
C14091 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__dfrtn_1_13/a_543_47# 0.00fF
C14092 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__inv_1_41/Y 0.01fF
C14093 sky130_fd_sc_hd__dfrtn_1_26/a_639_47# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C14094 sky130_fd_sc_hd__dfrtn_1_42/a_193_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C14095 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C14096 sky130_fd_sc_hd__nor3_2_3/C DOUT[15] 0.18fF
C14097 sky130_fd_sc_hd__dfrtn_1_27/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14098 sky130_fd_sc_hd__dfrtn_1_16/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14099 sky130_fd_sc_hd__dfrtn_1_8/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14100 sky130_fd_sc_hd__dfrtn_1_8/a_639_47# VDD 0.00fF
C14101 sky130_fd_sc_hd__dfrtn_1_3/a_1462_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C14102 sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# sky130_fd_sc_hd__inv_1_49/A 0.04fF
C14103 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C14104 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__nor3_1_19/a_193_297# 0.00fF
C14105 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__dfrtn_1_29/a_651_413# -0.00fF
C14106 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# sky130_fd_sc_hd__inv_1_7/A 0.01fF
C14107 DOUT[13] sky130_fd_sc_hd__dfrtn_1_34/a_761_289# 0.00fF
C14108 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__dfrtn_1_34/a_193_47# 0.00fF
C14109 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__dfrtn_1_34/a_27_47# 0.00fF
C14110 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# CLK_REF 0.01fF
C14111 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_20/a_1217_47# 0.00fF
C14112 sky130_fd_sc_hd__dfrtn_1_19/a_193_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C14113 sky130_fd_sc_hd__dfrtn_1_31/a_805_47# SEL_CONV_TIME[0] 0.00fF
C14114 sky130_fd_sc_hd__o311a_1_0/a_81_21# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C14115 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C14116 sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C14117 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14118 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__inv_1_44/A 0.02fF
C14119 sky130_fd_sc_hd__dfrtn_1_7/a_543_47# DOUT[14] 0.00fF
C14120 sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# sky130_fd_sc_hd__or3_1_0/C 0.01fF
C14121 sky130_fd_sc_hd__dfrtn_1_12/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14122 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__dfrtn_1_27/a_1270_413# 0.00fF
C14123 sky130_fd_sc_hd__nor3_2_0/a_27_297# VDD 0.06fF
C14124 sky130_fd_sc_hd__dfrtn_1_39/a_193_47# sky130_fd_sc_hd__inv_1_32/A 0.01fF
C14125 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__mux4_2_0/a_600_345# 0.01fF
C14126 sky130_fd_sc_hd__nor3_2_1/a_281_297# DOUT[15] 0.00fF
C14127 sky130_fd_sc_hd__dfrtn_1_7/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14128 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__inv_1_45/Y 0.15fF
C14129 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_3/a_639_47# 0.00fF
C14130 sky130_fd_sc_hd__dfrtn_1_7/a_1462_47# VDD 0.00fF
C14131 sky130_fd_sc_hd__dfrtn_1_17/a_448_47# RESET_COUNTERn 0.00fF
C14132 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# DOUT[14] 0.00fF
C14133 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__inv_1_54/A 0.01fF
C14134 sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C14135 DOUT[20] DOUT[14] 0.05fF
C14136 sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C14137 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_1108_47# 0.01fF
C14138 DOUT[4] sky130_fd_sc_hd__dfrtn_1_28/a_1217_47# 0.00fF
C14139 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__inv_1_7/A 0.01fF
C14140 sky130_fd_sc_hd__nor3_1_1/a_109_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14141 sky130_fd_sc_hd__inv_1_1/Y DOUT[18] 0.00fF
C14142 sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# sky130_fd_sc_hd__inv_1_0/Y 0.01fF
C14143 sky130_fd_sc_hd__nand3b_1_0/a_316_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C14144 DOUT[4] sky130_fd_sc_hd__dfrtn_1_35/a_27_47# 0.00fF
C14145 sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# sky130_fd_sc_hd__inv_1_11/Y 0.02fF
C14146 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# 0.00fF
C14147 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# 0.00fF
C14148 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_651_413# 0.00fF
C14149 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C14150 sky130_fd_sc_hd__mux4_2_0/a_1064_47# sky130_fd_sc_hd__nand2_1_1/Y 0.00fF
C14151 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__dfrtn_1_4/a_448_47# 0.00fF
C14152 DOUT[13] sky130_fd_sc_hd__inv_1_49/A 0.12fF
C14153 sky130_fd_sc_hd__dfrtn_1_31/a_1283_21# RESET_COUNTERn -0.00fF
C14154 sky130_fd_sc_hd__inv_1_37/A sky130_fd_sc_hd__inv_1_11/Y 0.01fF
C14155 sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C14156 sky130_fd_sc_hd__nor3_2_3/a_27_297# sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C14157 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C14158 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C14159 sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C14160 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14161 sky130_fd_sc_hd__or2_2_0/a_121_297# sky130_fd_sc_hd__dfrtn_1_19/a_543_47# 0.00fF
C14162 DOUT[11] VIN 0.20fF
C14163 sky130_fd_sc_hd__nor3_1_13/a_109_297# sky130_fd_sc_hd__dfrtn_1_10/a_448_47# 0.00fF
C14164 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C14165 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C14166 sky130_fd_sc_hd__dfrtn_1_11/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C14167 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C14168 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# sky130_fd_sc_hd__dfrtn_1_27/a_1462_47# 0.00fF
C14169 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# sky130_fd_sc_hd__dfrtn_1_27/a_1217_47# 0.00fF
C14170 sky130_fd_sc_hd__dfrtn_1_25/a_639_47# sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# 0.00fF
C14171 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_31/a_448_47# 0.00fF
C14172 sky130_fd_sc_hd__dfrtn_1_20/a_543_47# DOUT[2] 0.00fF
C14173 sky130_fd_sc_hd__o311a_1_0/a_585_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C14174 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__dfrtn_1_23/a_27_47# 0.00fF
C14175 sky130_fd_sc_hd__dfrtn_1_42/a_1462_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C14176 sky130_fd_sc_hd__dfrtn_1_31/a_761_289# DONE 0.00fF
C14177 sky130_fd_sc_hd__mux4_2_0/a_600_345# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C14178 sky130_fd_sc_hd__inv_1_37/A sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C14179 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# sky130_fd_sc_hd__inv_1_37/A 0.01fF
C14180 sky130_fd_sc_hd__nor3_1_12/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14181 sky130_fd_sc_hd__or3b_2_0/a_388_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14182 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# 0.01fF
C14183 sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C14184 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C14185 sky130_fd_sc_hd__dfrtn_1_23/a_805_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C14186 sky130_fd_sc_hd__dfrtn_1_32/a_639_47# RESET_COUNTERn 0.00fF
C14187 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__dfrtn_1_33/a_27_47# 0.00fF
C14188 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__dfrtn_1_33/a_448_47# 0.00fF
C14189 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__dfrtn_1_33/a_543_47# 0.00fF
C14190 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_33/a_761_289# 0.00fF
C14191 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_33/a_1108_47# 0.00fF
C14192 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__dfrtn_1_33/a_193_47# 0.00fF
C14193 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# SEL_CONV_TIME[0] 0.01fF
C14194 sky130_fd_sc_hd__o311a_1_0/a_266_297# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C14195 sky130_fd_sc_hd__dfrtn_1_31/a_639_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C14196 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# -0.00fF
C14197 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__dfrtn_1_14/a_448_47# -0.00fF
C14198 sky130_fd_sc_hd__dfrtn_1_28/a_651_413# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C14199 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__a221oi_4_0/a_1241_47# 0.00fF
C14200 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C14201 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# outb 0.00fF
C14202 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__dfrtn_1_22/a_805_47# -0.00fF
C14203 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# sky130_fd_sc_hd__dfrtn_1_22/a_639_47# -0.00fF
C14204 sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14205 sky130_fd_sc_hd__or3_1_0/C sky130_fd_sc_hd__inv_1_48/A 0.00fF
C14206 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# 0.00fF
C14207 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C14208 sky130_fd_sc_hd__dfrtn_1_24/a_1462_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C14209 sky130_fd_sc_hd__or2b_1_0/a_27_53# RESET_COUNTERn 0.00fF
C14210 sky130_fd_sc_hd__inv_1_38/Y RESET_COUNTERn 0.09fF
C14211 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C14212 sky130_fd_sc_hd__dfrtn_1_37/a_1270_413# VDD 0.00fF
C14213 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__inv_1_46/Y 0.00fF
C14214 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_17/a_639_47# 0.00fF
C14215 sky130_fd_sc_hd__or2b_1_0/X sky130_fd_sc_hd__inv_1_48/A 0.17fF
C14216 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__inv_1_11/Y 0.27fF
C14217 sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C14218 sky130_fd_sc_hd__dfrtn_1_3/a_651_413# VDD 0.01fF
C14219 sky130_fd_sc_hd__dfrtn_1_39/a_1462_47# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C14220 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# sky130_fd_sc_hd__inv_1_1/A 0.02fF
C14221 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C14222 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__dfrtp_1_2/a_193_47# 0.00fF
C14223 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__dfrtp_1_2/a_27_47# 0.00fF
C14224 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_2/a_543_47# 0.00fF
C14225 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_2/a_761_289# 0.00fF
C14226 sky130_fd_sc_hd__dfrtn_1_34/a_543_47# sky130_fd_sc_hd__inv_1_47/A 0.01fF
C14227 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C14228 sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__or2_2_0/X 0.00fF
C14229 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# RESET_COUNTERn 0.00fF
C14230 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_448_47# 0.00fF
C14231 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C14232 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C14233 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C14234 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C14235 sky130_fd_sc_hd__dfrtn_1_19/a_639_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C14236 DOUT[4] sky130_fd_sc_hd__dfrtn_1_35/a_1217_47# 0.00fF
C14237 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# DOUT[21] 0.00fF
C14238 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# 0.00fF
C14239 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_31/a_651_413# 0.00fF
C14240 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__dfrtn_1_23/a_193_47# -0.04fF
C14241 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__or3b_2_0/a_27_47# 0.00fF
C14242 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C14243 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# VDD 0.17fF
C14244 sky130_fd_sc_hd__dfrtn_1_9/a_543_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C14245 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14246 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.04fF
C14247 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# DOUT[11] 0.01fF
C14248 sky130_fd_sc_hd__dfrtn_1_4/a_543_47# VDD 0.05fF
C14249 sky130_fd_sc_hd__dfrtn_1_38/a_193_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C14250 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C14251 sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# 0.00fF
C14252 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# 0.00fF
C14253 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__dfrtn_1_26/a_651_413# 0.00fF
C14254 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# DOUT[3] 0.01fF
C14255 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C14256 sky130_fd_sc_hd__dfrtn_1_32/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14257 sky130_fd_sc_hd__dfrtn_1_25/a_805_47# SEL_CONV_TIME[1] 0.00fF
C14258 sky130_fd_sc_hd__dfrtn_1_21/a_805_47# VDD 0.00fF
C14259 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__or2_2_0/B 0.01fF
C14260 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C14261 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C14262 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_8/a_639_47# 0.00fF
C14263 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# 0.00fF
C14264 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# 0.00fF
C14265 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# 0.00fF
C14266 sky130_fd_sc_hd__dfrtn_1_19/a_448_47# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C14267 sky130_fd_sc_hd__inv_1_40/Y sky130_fd_sc_hd__inv_1_40/A 0.03fF
C14268 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_3/A 0.00fF
C14269 sky130_fd_sc_hd__dfrtn_1_16/a_193_47# sky130_fd_sc_hd__dfrtn_1_16/a_1108_47# -0.00fF
C14270 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# sky130_fd_sc_hd__dfrtn_1_16/a_448_47# -0.00fF
C14271 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C14272 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# DOUT[3] 0.00fF
C14273 sky130_fd_sc_hd__dfrtn_1_21/a_448_47# DOUT[2] 0.00fF
C14274 sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C14275 sky130_fd_sc_hd__dfrtn_1_38/a_805_47# sky130_fd_sc_hd__inv_1_27/Y 0.00fF
C14276 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# sky130_fd_sc_hd__o311a_1_0/A3 0.02fF
C14277 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C14278 DOUT[11] sky130_fd_sc_hd__inv_1_1/A 0.08fF
C14279 sky130_fd_sc_hd__inv_1_1/Y DOUT[22] 0.02fF
C14280 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C14281 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C14282 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_0/a_761_289# 0.04fF
C14283 sky130_fd_sc_hd__mux4_2_0/a_288_47# sky130_fd_sc_hd__inv_1_53/A 0.01fF
C14284 sky130_fd_sc_hd__dfrtn_1_28/a_193_47# sky130_fd_sc_hd__dfrtn_1_28/a_761_289# -0.00fF
C14285 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# sky130_fd_sc_hd__dfrtn_1_28/a_543_47# -0.00fF
C14286 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__dfrtn_1_16/a_1108_47# 0.00fF
C14287 sky130_fd_sc_hd__nor3_2_2/a_281_297# sky130_fd_sc_hd__dfrtn_1_16/a_1283_21# 0.00fF
C14288 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C14289 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__dfrtn_1_33/a_651_413# 0.00fF
C14290 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__dfrtn_1_33/a_1217_47# 0.00fF
C14291 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# VDD 0.11fF
C14292 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C14293 sky130_fd_sc_hd__dfrtp_1_3/a_639_47# RESET_COUNTERn 0.00fF
C14294 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_31/a_193_47# 0.00fF
C14295 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# -0.00fF
C14296 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# sky130_fd_sc_hd__dfrtn_1_6/a_543_47# -0.00fF
C14297 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__o211a_1_1/a_297_297# 0.00fF
C14298 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# RESET_COUNTERn 0.00fF
C14299 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C14300 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.00fF
C14301 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C14302 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.00fF
C14303 sky130_fd_sc_hd__dfrtn_1_39/a_761_289# VDD 0.06fF
C14304 sky130_fd_sc_hd__dfrtn_1_25/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14305 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14306 sky130_fd_sc_hd__dfrtn_1_25/a_639_47# VDD 0.00fF
C14307 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__nor3_2_0/a_27_297# 0.00fF
C14308 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_8/A 0.00fF
C14309 sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# sky130_fd_sc_hd__dfrtn_1_3/a_27_47# 0.00fF
C14310 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# 0.01fF
C14311 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__dfrtn_1_3/a_543_47# 0.00fF
C14312 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_3/a_651_413# 0.00fF
C14313 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__dfrtn_1_3/a_448_47# 0.00fF
C14314 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__dfrtn_1_3/a_193_47# 0.00fF
C14315 sky130_fd_sc_hd__dfrtn_1_41/a_448_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C14316 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C14317 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__nor3_2_3/C 0.44fF
C14318 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# sky130_fd_sc_hd__nor3_1_5/a_109_297# 0.00fF
C14319 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__nor3_1_5/a_193_297# 0.00fF
C14320 sky130_fd_sc_hd__o221ai_1_0/a_295_297# SEL_CONV_TIME[1] 0.00fF
C14321 sky130_fd_sc_hd__dfrtn_1_18/a_761_289# VDD 0.06fF
C14322 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__dfrtn_1_25/a_193_47# 0.00fF
C14323 sky130_fd_sc_hd__dfrtn_1_20/a_1270_413# sky130_fd_sc_hd__inv_1_35/Y 0.00fF
C14324 sky130_fd_sc_hd__inv_1_35/A DOUT[2] 0.03fF
C14325 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__inv_1_5/Y 0.03fF
C14326 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# DOUT[2] 0.00fF
C14327 VDD sky130_fd_sc_hd__inv_1_40/Y 0.51fF
C14328 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__dfrtp_1_2/a_651_413# 0.00fF
C14329 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C14330 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# 0.00fF
C14331 sky130_fd_sc_hd__dfrtn_1_24/a_651_413# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C14332 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__nor3_2_1/a_27_297# 0.00fF
C14333 sky130_fd_sc_hd__dfrtn_1_42/a_805_47# VDD -0.00fF
C14334 sky130_fd_sc_hd__dfrtn_1_42/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14335 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# DOUT[14] 0.01fF
C14336 sky130_fd_sc_hd__o311a_1_0/a_585_47# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C14337 sky130_fd_sc_hd__nor3_1_5/a_109_297# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C14338 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__nor3_1_4/a_193_297# 0.00fF
C14339 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_543_47# 0.00fF
C14340 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C14341 sky130_fd_sc_hd__dfrtn_1_29/a_805_47# RESET_COUNTERn 0.00fF
C14342 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C14343 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C14344 sky130_fd_sc_hd__dfrtn_1_38/a_193_47# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C14345 sky130_fd_sc_hd__dfrtn_1_10/a_639_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C14346 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C14347 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C14348 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# sky130_fd_sc_hd__dfrtn_1_38/a_543_47# 0.00fF
C14349 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_448_47# 0.00fF
C14350 sky130_fd_sc_hd__dfrtn_1_41/a_448_47# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C14351 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_36/a_805_47# 0.00fF
C14352 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__o311a_1_0/a_585_47# 0.00fF
C14353 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# DOUT[23] 0.00fF
C14354 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14355 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# VDD -0.00fF
C14356 sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14357 sky130_fd_sc_hd__nor3_1_3/a_109_297# RESET_COUNTERn 0.00fF
C14358 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_1/a_543_47# 0.00fF
C14359 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_1/a_193_47# 0.00fF
C14360 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# 0.00fF
C14361 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_805_47# 0.00fF
C14362 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__mux4_2_0/a_600_345# 0.00fF
C14363 sky130_fd_sc_hd__o311a_1_0/a_368_297# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C14364 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__nor3_2_3/C 0.33fF
C14365 sky130_fd_sc_hd__dfrtn_1_7/a_1462_47# DOUT[3] 0.00fF
C14366 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# 0.00fF
C14367 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C14368 sky130_fd_sc_hd__nor3_1_14/a_109_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14369 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# SEL_CONV_TIME[1] 0.02fF
C14370 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# sky130_fd_sc_hd__dfrtn_1_7/a_543_47# -0.00fF
C14371 sky130_fd_sc_hd__dfrtp_1_3/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14372 sky130_fd_sc_hd__dfrtn_1_16/a_448_47# DOUT[15] 0.01fF
C14373 sky130_fd_sc_hd__dfrtn_1_33/a_1108_47# sky130_fd_sc_hd__inv_1_43/A 0.01fF
C14374 sky130_fd_sc_hd__nor3_1_18/a_193_297# sky130_fd_sc_hd__inv_1_39/Y 0.00fF
C14375 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C14376 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C14377 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# RESET_COUNTERn 0.33fF
C14378 sky130_fd_sc_hd__dfrtn_1_26/a_543_47# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C14379 RESET_COUNTERn DOUT[18] 0.01fF
C14380 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__dfrtn_1_26/a_543_47# 0.00fF
C14381 sky130_fd_sc_hd__dfrtn_1_41/a_1270_413# sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C14382 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# sky130_fd_sc_hd__dfrtn_1_7/a_193_47# 0.00fF
C14383 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# sky130_fd_sc_hd__dfrtn_1_7/a_448_47# 0.00fF
C14384 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# sky130_fd_sc_hd__dfrtn_1_7/a_543_47# 0.00fF
C14385 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# 0.00fF
C14386 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_805_47# 0.00fF
C14387 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__dfrtn_1_7/a_651_413# 0.00fF
C14388 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# sky130_fd_sc_hd__dfrtn_1_7/a_27_47# 0.00fF
C14389 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__dfrtn_1_7/a_639_47# 0.00fF
C14390 DOUT[4] sky130_fd_sc_hd__dfrtn_1_12/a_448_47# 0.00fF
C14391 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__inv_1_0/Y 0.01fF
C14392 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# DOUT[20] 0.01fF
C14393 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# DOUT[6] 0.01fF
C14394 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C14395 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C14396 sky130_fd_sc_hd__nor3_1_5/A DOUT[4] 0.00fF
C14397 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__inv_1_0/Y 0.01fF
C14398 sky130_fd_sc_hd__dfrtp_1_0/a_1462_47# VDD 0.00fF
C14399 sky130_fd_sc_hd__dfrtp_1_0/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14400 sky130_fd_sc_hd__dfrtn_1_21/a_761_289# RESET_COUNTERn 0.02fF
C14401 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# DOUT[20] 0.00fF
C14402 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# RESET_COUNTERn 0.02fF
C14403 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# DOUT[8] 0.01fF
C14404 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# DOUT[7] 0.01fF
C14405 sky130_fd_sc_hd__dfrtn_1_22/a_1217_47# RESET_COUNTERn 0.00fF
C14406 sky130_fd_sc_hd__inv_1_11/Y DOUT[14] 0.00fF
C14407 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.00fF
C14408 VDD sky130_fd_sc_hd__inv_1_36/Y 0.35fF
C14409 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_32/a_448_47# 0.00fF
C14410 sky130_fd_sc_hd__o2111a_2_0/a_458_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C14411 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.00fF
C14412 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C14413 sky130_fd_sc_hd__dfrtn_1_30/a_1270_413# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C14414 sky130_fd_sc_hd__nor3_1_16/a_193_297# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C14415 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14416 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# VDD 0.06fF
C14417 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_10/a_639_47# -0.00fF
C14418 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.02fF
C14419 sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# outb 0.00fF
C14420 sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14421 sky130_fd_sc_hd__inv_1_30/A VDD 0.46fF
C14422 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__dfrtn_1_3/a_27_47# 0.00fF
C14423 sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C14424 sky130_fd_sc_hd__inv_1_37/A outb 0.02fF
C14425 sky130_fd_sc_hd__inv_1_3/Y DOUT[14] 0.01fF
C14426 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# DOUT[14] 0.01fF
C14427 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__inv_1_45/A 0.25fF
C14428 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C14429 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C14430 sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# sky130_fd_sc_hd__dfrtn_1_19/a_448_47# 0.00fF
C14431 sky130_fd_sc_hd__dfrtn_1_17/a_805_47# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C14432 sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# sky130_fd_sc_hd__inv_1_43/A 0.03fF
C14433 sky130_fd_sc_hd__dfrtn_1_16/a_639_47# RESET_COUNTERn 0.00fF
C14434 sky130_fd_sc_hd__inv_1_13/A sky130_fd_sc_hd__inv_1_5/A 0.19fF
C14435 sky130_fd_sc_hd__dfrtn_1_8/a_805_47# DOUT[21] 0.00fF
C14436 sky130_fd_sc_hd__dfrtn_1_8/a_1108_47# RESET_COUNTERn 0.01fF
C14437 CLK_REF sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C14438 sky130_fd_sc_hd__o311a_1_0/A3 DOUT[21] 0.01fF
C14439 sky130_fd_sc_hd__dfrtn_1_33/a_1462_47# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C14440 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__o211a_1_0/X 0.00fF
C14441 sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14442 sky130_fd_sc_hd__dfrtn_1_30/a_761_289# SEL_CONV_TIME[1] 0.01fF
C14443 VDD sky130_fd_sc_hd__dfrtn_1_9/a_805_47# 0.00fF
C14444 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_20/a_805_47# -0.00fF
C14445 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C14446 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# 0.00fF
C14447 sky130_fd_sc_hd__dfrtn_1_20/a_543_47# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C14448 sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C14449 sky130_fd_sc_hd__dfrtn_1_41/a_805_47# sky130_fd_sc_hd__dfrtn_1_38/a_651_413# 0.00fF
C14450 sky130_fd_sc_hd__dfrtn_1_41/a_651_413# sky130_fd_sc_hd__dfrtn_1_38/a_805_47# 0.00fF
C14451 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__dfrtn_1_38/a_1462_47# 0.00fF
C14452 sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C14453 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_13/a_543_47# 0.00fF
C14454 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_30/a_27_47# 0.00fF
C14455 sky130_fd_sc_hd__dfrtn_1_19/a_639_47# VDD 0.00fF
C14456 sky130_fd_sc_hd__dfrtp_1_3/a_1462_47# DOUT[23] 0.00fF
C14457 sky130_fd_sc_hd__nor3_1_0/a_109_297# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C14458 sky130_fd_sc_hd__dfrtn_1_26/a_543_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C14459 sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C14460 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C14461 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_18/a_639_47# 0.00fF
C14462 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C14463 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C14464 sky130_fd_sc_hd__dfrtn_1_31/a_448_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C14465 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_27/a_448_47# 0.00fF
C14466 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C14467 CLK_REF sky130_fd_sc_hd__or2_2_0/B 0.18fF
C14468 sky130_fd_sc_hd__dfrtn_1_23/a_1462_47# RESET_COUNTERn 0.00fF
C14469 sky130_fd_sc_hd__dfrtn_1_22/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14470 sky130_fd_sc_hd__nor3_1_3/a_109_297# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C14471 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__dfrtn_1_1/a_193_47# 0.00fF
C14472 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__inv_1_33/A 0.00fF
C14473 sky130_fd_sc_hd__dfrtn_1_7/a_805_47# DOUT[7] 0.00fF
C14474 sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# RESET_COUNTERn -0.00fF
C14475 sky130_fd_sc_hd__dfrtn_1_7/a_1462_47# DOUT[20] 0.00fF
C14476 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_29/a_651_413# 0.00fF
C14477 sky130_fd_sc_hd__dfrtn_1_10/a_1462_47# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C14478 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# DOUT[3] 0.00fF
C14479 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# VDD 0.10fF
C14480 sky130_fd_sc_hd__dfrtn_1_4/a_543_47# DOUT[3] 0.00fF
C14481 sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.00fF
C14482 sky130_fd_sc_hd__nor3_1_5/A outb 0.00fF
C14483 sky130_fd_sc_hd__dfrtn_1_16/a_193_47# DOUT[23] 0.00fF
C14484 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_27_47# 0.00fF
C14485 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_0/a_1217_47# -0.00fF
C14486 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# sky130_fd_sc_hd__dfrtn_1_0/a_805_47# -0.00fF
C14487 sky130_fd_sc_hd__dfrtn_1_14/a_761_289# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C14488 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__dfrtn_1_35/a_543_47# -0.00fF
C14489 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_2/A 0.01fF
C14490 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# CLK_REF 0.00fF
C14491 sky130_fd_sc_hd__dfrtn_1_4/a_543_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C14492 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# DOUT[17] 0.00fF
C14493 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_27_47# -0.00fF
C14494 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C14495 sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# sky130_fd_sc_hd__dfrtn_1_27/a_651_413# 0.00fF
C14496 sky130_fd_sc_hd__dfrtn_1_27/a_805_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C14497 sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C14498 sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.00fF
C14499 sky130_fd_sc_hd__nor3_2_2/a_27_297# DOUT[23] 0.00fF
C14500 sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14501 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C14502 sky130_fd_sc_hd__dfrtn_1_16/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14503 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14504 sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# VDD 0.00fF
C14505 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# SEL_CONV_TIME[0] 0.01fF
C14506 sky130_fd_sc_hd__dfrtn_1_8/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14507 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C14508 sky130_fd_sc_hd__dfrtn_1_36/a_543_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C14509 sky130_fd_sc_hd__dfrtn_1_17/a_193_47# sky130_fd_sc_hd__o211a_1_1/X 0.00fF
C14510 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C14511 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_31/a_1270_413# 0.00fF
C14512 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_27_47# 0.01fF
C14513 DOUT[22] RESET_COUNTERn 0.00fF
C14514 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C14515 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C14516 sky130_fd_sc_hd__nor3_1_17/a_109_297# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C14517 sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# DOUT[14] 0.00fF
C14518 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# 0.01fF
C14519 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__or2b_1_0/X 0.01fF
C14520 DOUT[4] sky130_fd_sc_hd__dfrtn_1_32/a_761_289# 0.00fF
C14521 VDD sky130_fd_sc_hd__o211a_1_1/X 0.58fF
C14522 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C14523 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__dfrtn_1_40/a_27_47# 0.00fF
C14524 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C14525 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# 0.00fF
C14526 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.01fF
C14527 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_17/a_543_47# 0.01fF
C14528 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__dfrtn_1_17/a_761_289# 0.00fF
C14529 sky130_fd_sc_hd__nor3_1_8/a_193_297# DOUT[14] 0.00fF
C14530 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# 0.00fF
C14531 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# 0.00fF
C14532 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__dfrtn_1_42/a_761_289# 0.00fF
C14533 sky130_fd_sc_hd__nor3_2_2/a_281_297# sky130_fd_sc_hd__dfrtn_1_42/a_193_47# 0.00fF
C14534 sky130_fd_sc_hd__dfrtn_1_20/a_448_47# sky130_fd_sc_hd__dfrtn_1_21/a_27_47# 0.00fF
C14535 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# sky130_fd_sc_hd__inv_1_6/A 0.01fF
C14536 sky130_fd_sc_hd__dfrtn_1_23/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14537 sky130_fd_sc_hd__nor3_1_13/a_193_297# VDD 0.00fF
C14538 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# 0.00fF
C14539 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__nor3_1_15/a_193_297# 0.00fF
C14540 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14541 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# VDD 0.10fF
C14542 sky130_fd_sc_hd__nor3_2_0/A DOUT[11] 0.00fF
C14543 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C14544 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# sky130_fd_sc_hd__o221ai_1_0/a_493_297# 0.00fF
C14545 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C14546 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C14547 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# sky130_fd_sc_hd__o221ai_1_0/a_295_297# 0.00fF
C14548 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.00fF
C14549 sky130_fd_sc_hd__dfrtn_1_7/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14550 sky130_fd_sc_hd__dfrtn_1_11/a_1217_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C14551 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# sky130_fd_sc_hd__inv_1_26/A 0.02fF
C14552 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__nor3_1_3/a_193_297# 0.00fF
C14553 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14554 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# VDD 0.00fF
C14555 sky130_fd_sc_hd__nor3_1_7/a_193_297# VIN 0.00fF
C14556 sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C14557 sky130_fd_sc_hd__dfrtn_1_42/a_1108_47# sky130_fd_sc_hd__dfrtn_1_23/a_193_47# 0.00fF
C14558 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_6/a_27_47# 0.01fF
C14559 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C14560 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# RESET_COUNTERn 0.00fF
C14561 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14562 sky130_fd_sc_hd__nor3_2_3/B DOUT[8] 0.02fF
C14563 sky130_fd_sc_hd__nor3_1_10/a_193_297# DOUT[8] 0.00fF
C14564 sky130_fd_sc_hd__nor3_1_10/a_109_297# RESET_COUNTERn 0.00fF
C14565 sky130_fd_sc_hd__dfrtn_1_33/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C14566 sky130_fd_sc_hd__dfrtn_1_33/a_651_413# VDD 0.00fF
C14567 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__nor3_1_19/Y 0.04fF
C14568 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# RESET_COUNTERn 0.02fF
C14569 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__nor3_1_4/A 0.01fF
C14570 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_5/Y 0.01fF
C14571 sky130_fd_sc_hd__dfrtn_1_22/a_448_47# sky130_fd_sc_hd__inv_1_40/Y 0.00fF
C14572 sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# VDD 0.00fF
C14573 sky130_fd_sc_hd__dfrtn_1_31/a_448_47# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C14574 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# DOUT[3] 0.00fF
C14575 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C14576 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__nor3_1_2/a_109_297# 0.00fF
C14577 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# VDD -0.16fF
C14578 sky130_fd_sc_hd__dfrtn_1_20/a_651_413# sky130_fd_sc_hd__inv_1_35/A 0.00fF
C14579 DOUT[4] sky130_fd_sc_hd__dfrtn_1_31/a_1270_413# 0.00fF
C14580 sky130_fd_sc_hd__inv_1_35/A sky130_fd_sc_hd__inv_1_30/Y 0.02fF
C14581 VDD DOUT[19] 1.22fF
C14582 sky130_fd_sc_hd__dfrtn_1_29/a_639_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C14583 sky130_fd_sc_hd__dfrtn_1_5/a_805_47# DOUT[14] 0.00fF
C14584 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C14585 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C14586 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__dfrtn_1_17/a_639_47# 0.00fF
C14587 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# HEADER_0/a_508_138# 0.00fF
C14588 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__or2_2_0/B 0.16fF
C14589 DOUT[13] DOUT[16] 0.03fF
C14590 DOUT[13] sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C14591 sky130_fd_sc_hd__dfrtn_1_0/a_761_289# DOUT[17] 0.00fF
C14592 sky130_fd_sc_hd__dfrtn_1_34/a_639_47# SEL_CONV_TIME[1] 0.00fF
C14593 sky130_fd_sc_hd__o211a_1_1/a_510_47# sky130_fd_sc_hd__dfrtn_1_17/a_651_413# 0.00fF
C14594 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__dfrtn_1_17/a_805_47# 0.00fF
C14595 sky130_fd_sc_hd__dfrtn_1_24/a_651_413# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C14596 sky130_fd_sc_hd__dfrtn_1_24/a_448_47# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C14597 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_651_413# 0.00fF
C14598 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_29/a_448_47# 0.00fF
C14599 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# DOUT[20] 0.01fF
C14600 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C14601 sky130_fd_sc_hd__nor3_1_5/a_109_297# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C14602 sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# VDD 0.07fF
C14603 sky130_fd_sc_hd__dfrtn_1_33/a_543_47# sky130_fd_sc_hd__inv_1_45/A 0.02fF
C14604 sky130_fd_sc_hd__inv_1_37/A sky130_fd_sc_hd__inv_1_13/Y 0.02fF
C14605 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_11/a_805_47# 0.00fF
C14606 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# 0.00fF
C14607 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__dfrtn_1_11/a_1270_413# 0.00fF
C14608 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# 0.00fF
C14609 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_1217_47# 0.00fF
C14610 sky130_fd_sc_hd__dfrtn_1_10/a_639_47# sky130_fd_sc_hd__dfrtn_1_11/a_761_289# 0.00fF
C14611 sky130_fd_sc_hd__nor3_2_3/a_281_297# VDD 0.04fF
C14612 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C14613 sky130_fd_sc_hd__dfrtn_1_42/a_543_47# DOUT[15] 0.00fF
C14614 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# 0.00fF
C14615 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/a_651_413# -0.00fF
C14616 sky130_fd_sc_hd__nor3_1_9/a_109_297# RESET_COUNTERn 0.00fF
C14617 sky130_fd_sc_hd__dfrtn_1_7/a_651_413# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C14618 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_17/a_1462_47# 0.00fF
C14619 sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# 0.00fF
C14620 sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# 0.00fF
C14621 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# 0.00fF
C14622 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__dfrtn_1_17/a_639_47# 0.00fF
C14623 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C14624 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_37/a_651_413# -0.00fF
C14625 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__dfrtn_1_37/a_448_47# -0.00fF
C14626 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_14/a_805_47# 0.00fF
C14627 sky130_fd_sc_hd__dfrtn_1_28/a_1270_413# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C14628 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14629 sky130_fd_sc_hd__inv_1_43/Y sky130_fd_sc_hd__nor3_2_3/B 0.04fF
C14630 sky130_fd_sc_hd__dfrtn_1_26/a_651_413# VDD 0.01fF
C14631 sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14632 sky130_fd_sc_hd__nor3_1_0/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14633 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# DOUT[14] 0.00fF
C14634 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__o2111a_2_0/X -0.03fF
C14635 sky130_fd_sc_hd__inv_1_6/A RESET_COUNTERn 0.46fF
C14636 sky130_fd_sc_hd__dfrtn_1_34/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14637 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C14638 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_41/a_193_47# -0.33fF
C14639 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C14640 sky130_fd_sc_hd__dfrtn_1_34/a_1270_413# VDD 0.00fF
C14641 sky130_fd_sc_hd__dfrtn_1_10/a_1462_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C14642 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# 0.00fF
C14643 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C14644 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_8/a_761_289# 0.01fF
C14645 sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C14646 sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# sky130_fd_sc_hd__inv_1_35/Y 0.01fF
C14647 sky130_fd_sc_hd__dfrtn_1_23/a_651_413# sky130_fd_sc_hd__inv_1_40/Y 0.01fF
C14648 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# -0.00fF
C14649 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# -0.00fF
C14650 sky130_fd_sc_hd__dfrtn_1_28/a_1270_413# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C14651 sky130_fd_sc_hd__dfrtn_1_41/a_651_413# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C14652 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__nand3b_1_0/Y 0.07fF
C14653 sky130_fd_sc_hd__inv_1_26/A DOUT[15] 0.40fF
C14654 sky130_fd_sc_hd__o221ai_1_0/a_493_297# SEL_CONV_TIME[0] 0.00fF
C14655 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__inv_1_50/A 0.26fF
C14656 sky130_fd_sc_hd__nor3_1_13/a_109_297# sky130_fd_sc_hd__inv_1_9/Y 0.00fF
C14657 sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# RESET_COUNTERn 0.01fF
C14658 sky130_fd_sc_hd__dfrtn_1_25/a_805_47# DOUT[21] 0.00fF
C14659 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C14660 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__or2_2_0/X 0.25fF
C14661 sky130_fd_sc_hd__inv_1_4/A DOUT[7] 0.00fF
C14662 sky130_fd_sc_hd__dfrtn_1_32/a_805_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C14663 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C14664 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__inv_1_32/Y 0.00fF
C14665 outb DOUT[14] 0.02fF
C14666 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C14667 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__o211a_1_1/a_215_47# 0.00fF
C14668 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__o211a_1_1/a_297_297# 0.00fF
C14669 VDD sky130_fd_sc_hd__inv_1_25/A 0.39fF
C14670 sky130_fd_sc_hd__dfrtp_1_0/a_1108_47# DOUT[15] 0.00fF
C14671 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C14672 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_26/a_543_47# 0.02fF
C14673 DOUT[13] sky130_fd_sc_hd__or3b_2_0/a_472_297# 0.00fF
C14674 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C14675 sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# HEADER_0/a_508_138# 0.00fF
C14676 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C14677 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C14678 sky130_fd_sc_hd__dfrtn_1_28/a_761_289# SEL_CONV_TIME[1] 0.00fF
C14679 sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# VDD 0.00fF
C14680 sky130_fd_sc_hd__dfrtn_1_42/a_448_47# RESET_COUNTERn 0.01fF
C14681 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# SEL_CONV_TIME[3] 0.01fF
C14682 sky130_fd_sc_hd__inv_1_52/Y sky130_fd_sc_hd__inv_1_36/A 0.01fF
C14683 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__o311a_1_0/a_266_47# 0.00fF
C14684 sky130_fd_sc_hd__dfrtn_1_34/a_805_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C14685 sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C14686 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_10/a_448_47# 0.01fF
C14687 sky130_fd_sc_hd__dfrtn_1_0/a_805_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C14688 sky130_fd_sc_hd__nor3_1_10/a_109_297# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C14689 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__or3_1_0/C 0.01fF
C14690 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtp_1_3/a_543_47# 0.00fF
C14691 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_651_413# 0.00fF
C14692 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__dfrtp_1_3/a_448_47# 0.00fF
C14693 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C14694 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C14695 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__mux4_2_0/a_788_316# -0.00fF
C14696 sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C14697 sky130_fd_sc_hd__o2111a_2_0/a_386_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14698 sky130_fd_sc_hd__o2111a_2_0/a_566_47# VDD 0.01fF
C14699 DOUT[13] sky130_fd_sc_hd__dfrtn_1_36/a_1462_47# 0.00fF
C14700 sky130_fd_sc_hd__nor3_1_20/a_193_297# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C14701 sky130_fd_sc_hd__nor3_1_4/A sky130_fd_sc_hd__inv_1_6/Y 0.17fF
C14702 sky130_fd_sc_hd__o221ai_1_0/a_213_123# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C14703 sky130_fd_sc_hd__dfrtn_1_17/a_805_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C14704 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# RESET_COUNTERn 0.00fF
C14705 sky130_fd_sc_hd__dfrtn_1_4/a_805_47# RESET_COUNTERn 0.00fF
C14706 sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# SEL_CONV_TIME[0] 0.00fF
C14707 sky130_fd_sc_hd__inv_1_49/Y SEL_CONV_TIME[0] 0.01fF
C14708 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_33/a_27_47# 0.00fF
C14709 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C14710 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__nor3_1_3/a_193_297# 0.00fF
C14711 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__nor3_1_3/a_109_297# 0.00fF
C14712 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14713 SLC_0/a_919_243# RESET_COUNTERn 0.06fF
C14714 sky130_fd_sc_hd__dfrtn_1_31/a_1108_47# sky130_fd_sc_hd__inv_1_49/A 0.03fF
C14715 DOUT[13] sky130_fd_sc_hd__dfrtn_1_31/a_543_47# 0.00fF
C14716 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_193_47# 0.00fF
C14717 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_27_47# 0.00fF
C14718 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# SEL_CONV_TIME[2] 0.02fF
C14719 SLC_0/a_438_293# lc_out 0.00fF
C14720 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_29/a_543_47# 0.01fF
C14721 sky130_fd_sc_hd__dfrtn_1_28/a_193_47# VDD 0.08fF
C14722 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C14723 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_761_289# -0.00fF
C14724 sky130_fd_sc_hd__dfrtn_1_14/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14725 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__nor3_1_13/a_193_297# 0.00fF
C14726 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C14727 sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# VDD 0.00fF
C14728 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# sky130_fd_sc_hd__dfrtn_1_0/a_1270_413# 0.00fF
C14729 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_0/a_1462_47# 0.00fF
C14730 sky130_fd_sc_hd__dfrtn_1_12/a_1270_413# sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# 0.00fF
C14731 sky130_fd_sc_hd__dfrtn_1_12/a_1462_47# sky130_fd_sc_hd__dfrtn_1_0/a_193_47# 0.00fF
C14732 sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C14733 CLK_REF sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# 0.00fF
C14734 sky130_fd_sc_hd__inv_1_23/A out 0.02fF
C14735 sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# DOUT[3] 0.00fF
C14736 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__dfrtn_1_29/a_761_289# 0.00fF
C14737 sky130_fd_sc_hd__dfrtp_1_0/a_1270_413# RESET_COUNTERn 0.00fF
C14738 sky130_fd_sc_hd__inv_1_15/A sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C14739 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_5/A 0.01fF
C14740 out RESET_COUNTERn 0.03fF
C14741 sky130_fd_sc_hd__o221ai_1_0/a_295_297# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C14742 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_38/a_1462_47# 0.00fF
C14743 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C14744 sky130_fd_sc_hd__inv_1_54/A RESET_COUNTERn 0.34fF
C14745 sky130_fd_sc_hd__dfrtn_1_3/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14746 sky130_fd_sc_hd__inv_1_48/A RESET_COUNTERn 1.05fF
C14747 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# lc_out 0.00fF
C14748 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C14749 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C14750 sky130_fd_sc_hd__inv_1_2/Y DOUT[6] 0.00fF
C14751 sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C14752 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__dfrtn_1_1/a_27_47# 0.00fF
C14753 sky130_fd_sc_hd__dfrtn_1_24/a_448_47# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C14754 sky130_fd_sc_hd__dfrtn_1_39/a_639_47# RESET_COUNTERn 0.00fF
C14755 sky130_fd_sc_hd__nor3_1_14/a_109_297# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C14756 sky130_fd_sc_hd__dfrtn_1_22/a_651_413# sky130_fd_sc_hd__inv_1_39/Y 0.00fF
C14757 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__inv_1_13/A 0.04fF
C14758 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# DOUT[21] 0.01fF
C14759 sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C14760 sky130_fd_sc_hd__o311a_1_0/a_81_21# sky130_fd_sc_hd__nand2_1_1/a_113_47# 0.00fF
C14761 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__inv_1_42/A 0.02fF
C14762 sky130_fd_sc_hd__dfrtp_1_3/a_1462_47# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C14763 sky130_fd_sc_hd__nor3_1_16/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14764 sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C14765 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__o2111a_2_0/a_80_21# 0.00fF
C14766 sky130_fd_sc_hd__dfrtn_1_18/a_639_47# RESET_COUNTERn 0.00fF
C14767 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C14768 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__inv_1_6/A 0.01fF
C14769 DONE sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C14770 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__dfrtn_1_25/a_543_47# 0.00fF
C14771 sky130_fd_sc_hd__or3_1_0/a_111_297# sky130_fd_sc_hd__dfrtn_1_25/a_761_289# 0.00fF
C14772 sky130_fd_sc_hd__or3_1_0/a_183_297# sky130_fd_sc_hd__dfrtn_1_25/a_193_47# 0.00fF
C14773 sky130_fd_sc_hd__dfrtn_1_20/a_761_289# sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# 0.00fF
C14774 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C14775 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C14776 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C14777 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C14778 sky130_fd_sc_hd__dfrtn_1_4/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14779 DOUT[4] SEL_CONV_TIME[0] 0.53fF
C14780 sky130_fd_sc_hd__dfrtn_1_30/a_543_47# SEL_CONV_TIME[0] 0.02fF
C14781 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# 0.00fF
C14782 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# 0.00fF
C14783 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__dfrtn_1_7/a_193_47# 0.00fF
C14784 sky130_fd_sc_hd__mux4_1_0/a_27_413# VDD 0.03fF
C14785 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# DOUT[3] 0.00fF
C14786 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__nor3_1_4/A 0.01fF
C14787 SLC_0/a_438_293# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C14788 sky130_fd_sc_hd__dfrtn_1_10/a_1283_21# VDD 0.11fF
C14789 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14790 sky130_fd_sc_hd__dfrtn_1_9/a_448_47# RESET_COUNTERn 0.00fF
C14791 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_761_289# 0.00fF
C14792 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_193_47# 0.00fF
C14793 sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# sky130_fd_sc_hd__dfrtp_1_3/a_651_413# 0.00fF
C14794 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# DOUT[23] 0.00fF
C14795 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__mux4_2_0/a_1064_47# -0.00fF
C14796 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C14797 sky130_fd_sc_hd__dfrtn_1_19/a_1108_47# RESET_COUNTERn 0.00fF
C14798 CLK_REF sky130_fd_sc_hd__dfrtn_1_17/a_639_47# 0.00fF
C14799 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C14800 sky130_fd_sc_hd__o311a_1_0/a_368_297# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C14801 sky130_fd_sc_hd__mux4_2_0/a_193_47# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C14802 sky130_fd_sc_hd__nor3_1_17/a_193_297# RESET_COUNTERn 0.00fF
C14803 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C14804 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_761_289# -0.00fF
C14805 sky130_fd_sc_hd__mux4_2_0/a_193_369# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C14806 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14807 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__dfrtn_1_4/a_761_289# 0.00fF
C14808 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_4/a_543_47# 0.00fF
C14809 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C14810 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.01fF
C14811 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__inv_1_8/A 0.02fF
C14812 sky130_fd_sc_hd__dfrtn_1_21/a_1462_47# RESET_COUNTERn 0.00fF
C14813 sky130_fd_sc_hd__inv_1_50/Y sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14814 sky130_fd_sc_hd__dfrtn_1_35/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_1270_413# 0.00fF
C14815 sky130_fd_sc_hd__dfrtn_1_35/a_448_47# sky130_fd_sc_hd__dfrtn_1_36/a_543_47# 0.00fF
C14816 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_639_47# 0.00fF
C14817 DOUT[19] DOUT[3] 0.04fF
C14818 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# 0.00fF
C14819 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_1217_47# 0.00fF
C14820 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# 0.00fF
C14821 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_1462_47# 0.00fF
C14822 sky130_fd_sc_hd__nor3_1_2/a_109_297# RESET_COUNTERn 0.00fF
C14823 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C14824 sky130_fd_sc_hd__dfrtn_1_28/a_1462_47# VDD 0.00fF
C14825 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C14826 sky130_fd_sc_hd__inv_1_47/Y SEL_CONV_TIME[0] 0.19fF
C14827 sky130_fd_sc_hd__dfrtn_1_27/a_761_289# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C14828 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_37/a_651_413# 0.00fF
C14829 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C14830 sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C14831 sky130_fd_sc_hd__dfrtn_1_21/a_1217_47# DOUT[2] 0.00fF
C14832 sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# VDD 0.08fF
C14833 sky130_fd_sc_hd__dfrtn_1_0/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C14834 sky130_fd_sc_hd__dfrtn_1_35/a_193_47# VDD 0.10fF
C14835 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__inv_1_15/A 0.24fF
C14836 sky130_fd_sc_hd__inv_1_2/A DOUT[19] 0.04fF
C14837 sky130_fd_sc_hd__nor3_1_13/a_193_297# sky130_fd_sc_hd__dfrtn_1_8/a_27_47# 0.00fF
C14838 sky130_fd_sc_hd__nor3_1_13/a_109_297# sky130_fd_sc_hd__dfrtn_1_8/a_193_47# 0.00fF
C14839 sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# sky130_fd_sc_hd__inv_1_14/A 0.02fF
C14840 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# DOUT[17] 0.00fF
C14841 sky130_fd_sc_hd__nor3_1_3/a_109_297# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C14842 sky130_fd_sc_hd__mux4_1_0/a_834_97# SEL_CONV_TIME[1] 0.00fF
C14843 sky130_fd_sc_hd__nor3_2_0/A sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C14844 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_38/a_639_47# 0.00fF
C14845 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C14846 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# sky130_fd_sc_hd__or3_1_0/C 0.53fF
C14847 HEADER_0/a_508_138# sky130_fd_sc_hd__inv_1_6/A 0.01fF
C14848 sky130_fd_sc_hd__nor3_1_5/a_193_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14849 sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C14850 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# 0.00fF
C14851 sky130_fd_sc_hd__dfrtn_1_23/a_761_289# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C14852 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C14853 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_24/a_193_47# 0.00fF
C14854 sky130_fd_sc_hd__dfrtn_1_39/a_448_47# sky130_fd_sc_hd__inv_1_32/Y -0.02fF
C14855 sky130_fd_sc_hd__dfrtn_1_20/a_805_47# VDD 0.00fF
C14856 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# RESET_COUNTERn 0.00fF
C14857 sky130_fd_sc_hd__inv_1_13/Y DOUT[14] 0.36fF
C14858 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_761_289# -0.00fF
C14859 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# RESET_COUNTERn 0.02fF
C14860 sky130_fd_sc_hd__dfrtn_1_25/a_1462_47# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C14861 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C14862 sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14863 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# SEL_CONV_TIME[1] 0.00fF
C14864 CLK_REF sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.04fF
C14865 sky130_fd_sc_hd__inv_1_48/A SEL_CONV_TIME[3] 0.01fF
C14866 DOUT[1] sky130_fd_sc_hd__dfrtn_1_36/a_805_47# 0.00fF
C14867 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# 0.03fF
C14868 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_4/a_651_413# 0.00fF
C14869 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__inv_1_31/A 0.00fF
C14870 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# -0.00fF
C14871 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_12/a_543_47# -0.00fF
C14872 sky130_fd_sc_hd__dfrtn_1_16/a_651_413# DOUT[2] 0.00fF
C14873 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# 0.00fF
C14874 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__dfrtn_1_13/a_761_289# 0.00fF
C14875 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# 0.00fF
C14876 DOUT[9] sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C14877 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# sky130_fd_sc_hd__dfrtn_1_42/a_1217_47# -0.00fF
C14878 DOUT[9] sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.01fF
C14879 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# DOUT[11] 0.00fF
C14880 sky130_fd_sc_hd__nor3_1_18/a_193_297# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C14881 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__dfrtp_1_0/a_543_47# -0.00fF
C14882 DOUT[1] sky130_fd_sc_hd__nor3_2_3/C 0.51fF
C14883 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14884 sky130_fd_sc_hd__mux4_1_0/a_668_97# VDD 0.00fF
C14885 sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__nor3_2_3/C 0.13fF
C14886 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C14887 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C14888 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C14889 sky130_fd_sc_hd__o211a_1_0/a_215_47# sky130_fd_sc_hd__nor3_2_3/C 0.03fF
C14890 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# VIN 0.03fF
C14891 sky130_fd_sc_hd__dfrtp_1_0/a_1217_47# DOUT[23] 0.00fF
C14892 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C14893 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__inv_1_51/Y 0.07fF
C14894 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C14895 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_639_47# -0.00fF
C14896 sky130_fd_sc_hd__or2_2_0/a_121_297# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C14897 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C14898 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# RESET_COUNTERn 0.00fF
C14899 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_11/a_1270_413# 0.00fF
C14900 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C14901 SEL_CONV_TIME[2] sky130_fd_sc_hd__inv_1_48/A 0.00fF
C14902 sky130_fd_sc_hd__dfrtn_1_38/a_651_413# SEL_CONV_TIME[0] 0.00fF
C14903 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# VDD 0.23fF
C14904 sky130_fd_sc_hd__nor3_2_0/a_27_297# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C14905 sky130_fd_sc_hd__mux4_2_0/a_1281_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C14906 sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C14907 DOUT[4] sky130_fd_sc_hd__nor3_2_0/a_27_297# 0.00fF
C14908 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# RESET_COUNTERn 0.00fF
C14909 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# DOUT[20] 0.00fF
C14910 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# sky130_fd_sc_hd__dfrtn_1_4/a_448_47# 0.00fF
C14911 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_448_47# -0.00fF
C14912 sky130_fd_sc_hd__dfrtn_1_39/a_639_47# SEL_CONV_TIME[2] 0.00fF
C14913 sky130_fd_sc_hd__nor3_1_19/Y sky130_fd_sc_hd__inv_1_44/A 0.06fF
C14914 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C14915 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_39/a_193_47# 0.00fF
C14916 sky130_fd_sc_hd__or2b_1_0/X sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C14917 sky130_fd_sc_hd__or2_2_0/B sky130_fd_sc_hd__nor3_2_3/C 0.06fF
C14918 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__o311a_1_0/a_585_47# 0.00fF
C14919 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__inv_1_45/A 0.00fF
C14920 sky130_fd_sc_hd__dfrtn_1_39/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# 0.00fF
C14921 sky130_fd_sc_hd__dfrtn_1_33/a_543_47# RESET_COUNTERn 0.00fF
C14922 DOUT[1] sky130_fd_sc_hd__dfrtn_1_32/a_448_47# 0.00fF
C14923 sky130_fd_sc_hd__dfrtn_1_7/a_543_47# DOUT[19] 0.00fF
C14924 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__dfrtn_1_14/a_193_47# 0.00fF
C14925 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__dfrtn_1_14/a_27_47# 0.00fF
C14926 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C14927 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_30/a_27_47# 0.01fF
C14928 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C14929 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__mux4_2_0/a_872_316# 0.00fF
C14930 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__mux4_2_0/a_600_345# 0.00fF
C14931 sky130_fd_sc_hd__dfrtn_1_35/a_1462_47# VDD 0.00fF
C14932 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__inv_1_34/A 0.00fF
C14933 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C14934 sky130_fd_sc_hd__dfrtn_1_30/a_1270_413# RESET_COUNTERn 0.00fF
C14935 sky130_fd_sc_hd__dfrtn_1_12/a_1462_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C14936 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.00fF
C14937 SLC_0/a_264_22# SLC_0/a_919_243# -0.00fF
C14938 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__inv_1_8/Y 0.03fF
C14939 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C14940 sky130_fd_sc_hd__dfrtn_1_3/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.00fF
C14941 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C14942 sky130_fd_sc_hd__nor3_1_11/a_193_297# VDD 0.00fF
C14943 sky130_fd_sc_hd__dfrtn_1_18/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# -0.00fF
C14944 sky130_fd_sc_hd__dfrtn_1_18/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_448_47# -0.00fF
C14945 sky130_fd_sc_hd__mux4_2_0/a_1060_369# SEL_CONV_TIME[1] 0.00fF
C14946 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# DOUT[19] 0.00fF
C14947 sky130_fd_sc_hd__dfrtn_1_27/a_1217_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C14948 DOUT[19] DOUT[20] 0.03fF
C14949 sky130_fd_sc_hd__dfrtn_1_34/a_805_47# SEL_CONV_TIME[0] 0.00fF
C14950 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C14951 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__inv_1_34/Y 0.01fF
C14952 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14953 sky130_fd_sc_hd__dfrtp_1_1/a_639_47# VDD 0.00fF
C14954 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__inv_1_31/Y 0.14fF
C14955 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_30/a_805_47# 0.00fF
C14956 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C14957 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__nor3_1_0/A 0.19fF
C14958 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C14959 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C14960 sky130_fd_sc_hd__dfrtn_1_30/a_448_47# DONE 0.00fF
C14961 sky130_fd_sc_hd__dfrtn_1_16/a_1283_21# sky130_fd_sc_hd__inv_1_25/A 0.01fF
C14962 sky130_fd_sc_hd__dfrtp_1_0/a_1270_413# SLC_0/a_264_22# 0.00fF
C14963 sky130_fd_sc_hd__dfrtp_1_0/a_639_47# SLC_0/a_438_293# 0.00fF
C14964 sky130_fd_sc_hd__inv_1_38/A sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C14965 SLC_0/a_264_22# out 0.02fF
C14966 sky130_fd_sc_hd__dfrtn_1_38/a_193_47# RESET_COUNTERn 0.29fF
C14967 sky130_fd_sc_hd__dfrtn_1_14/a_543_47# DOUT[18] 0.00fF
C14968 sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# SEL_CONV_TIME[1] 0.00fF
C14969 sky130_fd_sc_hd__dfrtn_1_42/a_1462_47# sky130_fd_sc_hd__inv_1_40/Y 0.00fF
C14970 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C14971 CLK_REF sky130_fd_sc_hd__dfrtp_1_3/a_1462_47# 0.00fF
C14972 sky130_fd_sc_hd__nor3_2_1/a_281_297# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C14973 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# 0.00fF
C14974 sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# sky130_fd_sc_hd__or2_2_0/a_121_297# 0.00fF
C14975 sky130_fd_sc_hd__dfrtn_1_8/a_639_47# outb 0.00fF
C14976 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_10/a_1283_21# 0.02fF
C14977 DOUT[9] sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# 0.00fF
C14978 sky130_fd_sc_hd__dfrtn_1_39/a_193_47# sky130_fd_sc_hd__inv_1_33/A 0.02fF
C14979 sky130_fd_sc_hd__dfrtn_1_7/a_805_47# VIN 0.00fF
C14980 sky130_fd_sc_hd__o311a_1_0/a_585_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14981 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_14/A 0.01fF
C14982 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_12/a_639_47# 0.00fF
C14983 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C14984 sky130_fd_sc_hd__mux4_2_0/a_600_345# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C14985 sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# DOUT[5] 0.00fF
C14986 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C14987 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C14988 sky130_fd_sc_hd__mux4_2_0/a_872_316# VDD 0.03fF
C14989 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# out 0.00fF
C14990 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_21/a_193_47# 0.00fF
C14991 sky130_fd_sc_hd__dfrtn_1_18/a_193_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C14992 sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# SEL_CONV_TIME[1] 0.00fF
C14993 sky130_fd_sc_hd__dfrtn_1_26/a_543_47# RESET_COUNTERn 0.02fF
C14994 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_2/a_543_47# 0.02fF
C14995 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# sky130_fd_sc_hd__inv_1_53/A 0.02fF
C14996 sky130_fd_sc_hd__dfrtn_1_34/a_1462_47# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C14997 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C14998 sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C14999 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C15000 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_3/a_761_289# 0.00fF
C15001 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C15002 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C15003 sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C15004 sky130_fd_sc_hd__dfrtn_1_35/a_651_413# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C15005 sky130_fd_sc_hd__dfrtn_1_16/a_761_289# sky130_fd_sc_hd__nor3_2_3/A 0.02fF
C15006 sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15007 sky130_fd_sc_hd__dfrtn_1_34/a_639_47# DOUT[21] 0.00fF
C15008 sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# RESET_COUNTERn 0.03fF
C15009 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15010 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# VDD 0.01fF
C15011 sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# RESET_COUNTERn 0.00fF
C15012 sky130_fd_sc_hd__dfrtn_1_35/a_448_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C15013 sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# VDD 0.00fF
C15014 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C15015 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C15016 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# DOUT[2] 0.00fF
C15017 sky130_fd_sc_hd__nor3_2_0/a_27_297# outb 0.00fF
C15018 sky130_fd_sc_hd__nor3_2_2/a_281_297# sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C15019 sky130_fd_sc_hd__dfrtn_1_8/a_1283_21# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C15020 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_35/a_193_47# 0.00fF
C15021 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_39/a_1462_47# 0.00fF
C15022 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# DONE 0.00fF
C15023 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# 0.00fF
C15024 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__nand3b_1_0/a_53_93# 0.01fF
C15025 sky130_fd_sc_hd__mux4_2_0/a_1279_413# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C15026 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C15027 sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# VDD 0.10fF
C15028 sky130_fd_sc_hd__dfrtn_1_27/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15029 sky130_fd_sc_hd__dfrtp_1_3/a_448_47# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C15030 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# 0.00fF
C15031 sky130_fd_sc_hd__dfrtn_1_34/a_639_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C15032 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C15033 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# RESET_COUNTERn 0.01fF
C15034 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__dfrtn_1_1/a_543_47# 0.00fF
C15035 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__dfrtn_1_1/a_761_289# 0.00fF
C15036 sky130_fd_sc_hd__o211a_1_1/a_510_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15037 sky130_fd_sc_hd__dfrtn_1_37/a_1462_47# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C15038 sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C15039 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# -0.00fF
C15040 sky130_fd_sc_hd__dfrtn_1_36/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_543_47# -0.00fF
C15041 sky130_fd_sc_hd__inv_1_36/A sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15042 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C15043 sky130_fd_sc_hd__dfrtn_1_29/a_805_47# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C15044 sky130_fd_sc_hd__o2111a_2_0/a_80_21# RESET_COUNTERn 0.00fF
C15045 sky130_fd_sc_hd__nor3_1_3/a_193_297# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C15046 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C15047 sky130_fd_sc_hd__dfrtn_1_38/a_1462_47# RESET_COUNTERn 0.00fF
C15048 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# sky130_fd_sc_hd__inv_1_43/Y 0.02fF
C15049 sky130_fd_sc_hd__nor3_1_10/a_109_297# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C15050 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__or3b_2_0/X 0.02fF
C15051 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# DOUT[18] 0.00fF
C15052 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C15053 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C15054 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# VDD 0.01fF
C15055 DOUT[13] RESET_COUNTERn 0.10fF
C15056 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.00fF
C15057 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_639_47# 0.00fF
C15058 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C15059 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_805_47# 0.00fF
C15060 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C15061 sky130_fd_sc_hd__dfrtp_1_3/a_448_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C15062 sky130_fd_sc_hd__nor3_1_15/a_193_297# DOUT[1] 0.00fF
C15063 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__nor3_1_1/a_109_297# 0.00fF
C15064 sky130_fd_sc_hd__a221oi_4_0/a_27_297# SEL_CONV_TIME[1] 0.00fF
C15065 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C15066 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.01fF
C15067 sky130_fd_sc_hd__dfrtn_1_12/a_651_413# VDD 0.01fF
C15068 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15069 sky130_fd_sc_hd__inv_1_41/Y sky130_fd_sc_hd__nor3_2_3/B 0.16fF
C15070 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C15071 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# 0.00fF
C15072 sky130_fd_sc_hd__dfrtp_1_2/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15073 sky130_fd_sc_hd__dfrtn_1_39/a_1462_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C15074 sky130_fd_sc_hd__dfrtn_1_17/a_1270_413# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C15075 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_1/a_193_47# 0.00fF
C15076 sky130_fd_sc_hd__inv_1_8/A RESET_COUNTERn 1.47fF
C15077 sky130_fd_sc_hd__dfrtn_1_28/a_761_289# DOUT[21] 0.00fF
C15078 sky130_fd_sc_hd__dfrtn_1_33/a_448_47# DOUT[23] 0.00fF
C15079 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__nor3_1_1/a_193_297# 0.00fF
C15080 sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# DOUT[5] 0.00fF
C15081 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# -0.00fF
C15082 sky130_fd_sc_hd__mux4_1_0/a_247_21# SEL_CONV_TIME[0] 0.00fF
C15083 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# RESET_COUNTERn 0.01fF
C15084 sky130_fd_sc_hd__or3_1_0/X sky130_fd_sc_hd__inv_1_48/A 0.18fF
C15085 DONE sky130_fd_sc_hd__inv_1_49/A 0.18fF
C15086 sky130_fd_sc_hd__dfrtn_1_28/a_448_47# sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C15087 sky130_fd_sc_hd__dfrtn_1_18/a_1462_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C15088 sky130_fd_sc_hd__dfrtn_1_42/a_448_47# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C15089 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_34/a_651_413# 0.00fF
C15090 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C15091 sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C15092 sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# sky130_fd_sc_hd__dfrtp_1_3/a_761_289# 0.00fF
C15093 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__dfrtp_1_3/a_448_47# 0.00fF
C15094 sky130_fd_sc_hd__dfrtp_1_1/a_639_47# sky130_fd_sc_hd__o211a_1_0/X 0.00fF
C15095 sky130_fd_sc_hd__dfrtn_1_33/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15096 sky130_fd_sc_hd__dfrtn_1_21/a_1217_47# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C15097 sky130_fd_sc_hd__dfrtn_1_20/a_651_413# sky130_fd_sc_hd__dfrtn_1_21/a_1217_47# 0.00fF
C15098 sky130_fd_sc_hd__dfrtn_1_36/a_651_413# sky130_fd_sc_hd__inv_1_40/A 0.00fF
C15099 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__nand3b_1_1/a_316_47# 0.00fF
C15100 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# VIN 0.00fF
C15101 sky130_fd_sc_hd__dfrtn_1_14/a_543_47# DOUT[22] 0.00fF
C15102 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__dfrtn_1_34/a_27_47# 0.00fF
C15103 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__dfrtn_1_34/a_193_47# 0.00fF
C15104 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# 0.00fF
C15105 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_37/a_543_47# 0.00fF
C15106 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# sky130_fd_sc_hd__dfrtn_1_37/a_193_47# 0.00fF
C15107 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# sky130_fd_sc_hd__dfrtn_1_37/a_27_47# 0.00fF
C15108 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_37/a_651_413# 0.00fF
C15109 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_37/a_639_47# 0.00fF
C15110 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_37/a_805_47# 0.00fF
C15111 sky130_fd_sc_hd__dfrtn_1_40/a_1270_413# sky130_fd_sc_hd__dfrtn_1_37/a_761_289# 0.00fF
C15112 sky130_fd_sc_hd__nor3_1_1/a_109_297# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C15113 sky130_fd_sc_hd__inv_1_46/Y DOUT[23] 0.00fF
C15114 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15115 sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C15116 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C15117 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C15118 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_805_47# 0.00fF
C15119 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_2/a_651_413# 0.00fF
C15120 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_639_47# 0.00fF
C15121 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__dfrtn_1_2/a_448_47# 0.00fF
C15122 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__dfrtn_1_2/a_543_47# 0.00fF
C15123 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# 0.00fF
C15124 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_25/a_193_47# 0.00fF
C15125 sky130_fd_sc_hd__dfrtn_1_22/a_761_289# sky130_fd_sc_hd__inv_1_39/A 0.01fF
C15126 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_24/a_448_47# -0.00fF
C15127 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# -0.00fF
C15128 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# 0.00fF
C15129 VDD SEL_CONV_TIME[1] 3.23fF
C15130 sky130_fd_sc_hd__dfrtn_1_38/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15131 sky130_fd_sc_hd__inv_1_4/Y sky130_fd_sc_hd__inv_1_6/A 0.11fF
C15132 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__inv_1_49/A 0.39fF
C15133 DOUT[1] sky130_fd_sc_hd__dfrtn_1_22/a_1270_413# 0.00fF
C15134 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_34/a_193_47# 0.01fF
C15135 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# -0.03fF
C15136 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# RESET_COUNTERn 0.03fF
C15137 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# 0.02fF
C15138 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.02fF
C15139 sky130_fd_sc_hd__dfrtn_1_26/a_448_47# DOUT[23] 0.00fF
C15140 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# DOUT[14] 0.00fF
C15141 sky130_fd_sc_hd__inv_1_24/A sky130_fd_sc_hd__inv_1_23/A 0.18fF
C15142 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# DOUT[19] 0.01fF
C15143 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__inv_1_15/A 0.01fF
C15144 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# 0.00fF
C15145 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__dfrtn_1_15/a_193_47# 0.00fF
C15146 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C15147 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__dfrtn_1_15/a_27_47# 0.00fF
C15148 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_651_413# 0.00fF
C15149 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# 0.00fF
C15150 sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C15151 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C15152 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# 0.00fF
C15153 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C15154 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C15155 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C15156 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_639_47# 0.00fF
C15157 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C15158 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C15159 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# VDD 0.17fF
C15160 sky130_fd_sc_hd__dfrtn_1_3/a_761_289# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C15161 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# sky130_fd_sc_hd__nor3_1_0/a_193_297# 0.00fF
C15162 sky130_fd_sc_hd__dfrtn_1_14/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C15163 sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15164 sky130_fd_sc_hd__dfrtn_1_36/a_651_413# VDD 0.01fF
C15165 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# 0.00fF
C15166 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# 0.00fF
C15167 sky130_fd_sc_hd__inv_1_4/A VIN 0.03fF
C15168 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__nor3_1_19/Y 0.01fF
C15169 sky130_fd_sc_hd__or2b_1_0/a_301_297# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C15170 sky130_fd_sc_hd__nor3_2_3/a_281_297# sky130_fd_sc_hd__dfrtn_1_42/a_193_47# 0.00fF
C15171 sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15172 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_13/a_761_289# 0.00fF
C15173 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C15174 sky130_fd_sc_hd__dfrtn_1_17/a_651_413# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C15175 sky130_fd_sc_hd__dfrtn_1_0/a_639_47# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C15176 sky130_fd_sc_hd__nor3_1_13/a_193_297# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C15177 sky130_fd_sc_hd__nor3_1_11/a_193_297# DOUT[3] 0.00fF
C15178 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C15179 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__inv_1_53/A 0.00fF
C15180 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C15181 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C15182 SEL_CONV_TIME[0] sky130_fd_sc_hd__inv_1_44/A 0.29fF
C15183 sky130_fd_sc_hd__o2111a_2_0/a_80_21# SEL_CONV_TIME[3] 0.01fF
C15184 sky130_fd_sc_hd__dfrtn_1_28/a_1270_413# RESET_COUNTERn -0.00fF
C15185 sky130_fd_sc_hd__dfrtn_1_39/a_639_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C15186 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C15187 sky130_fd_sc_hd__dfrtn_1_30/a_639_47# sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C15188 sky130_fd_sc_hd__nor3_1_11/a_193_297# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C15189 sky130_fd_sc_hd__nor3_1_3/a_193_297# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C15190 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# RESET_COUNTERn 0.00fF
C15191 sky130_fd_sc_hd__dfrtn_1_35/a_761_289# DOUT[21] 0.00fF
C15192 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__inv_1_41/Y 0.19fF
C15193 sky130_fd_sc_hd__inv_1_29/Y sky130_fd_sc_hd__o211a_1_1/X 0.08fF
C15194 DOUT[4] sky130_fd_sc_hd__inv_1_36/Y 0.44fF
C15195 sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C15196 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__or2b_1_0/X 0.01fF
C15197 sky130_fd_sc_hd__dfrtn_1_23/a_543_47# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C15198 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C15199 sky130_fd_sc_hd__inv_1_27/Y RESET_COUNTERn 0.02fF
C15200 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_39/a_193_47# 0.00fF
C15201 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# 0.00fF
C15202 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_543_47# 0.00fF
C15203 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# SEL_CONV_TIME[2] 0.00fF
C15204 sky130_fd_sc_hd__conb_1_0/LO sky130_fd_sc_hd__nor3_2_3/B 0.03fF
C15205 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_30/a_193_47# 0.01fF
C15206 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C15207 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# 0.00fF
C15208 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C15209 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C15210 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_448_47# 0.00fF
C15211 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C15212 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_761_289# 0.00fF
C15213 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C15214 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# DOUT[22] 0.00fF
C15215 sky130_fd_sc_hd__dfrtn_1_20/a_448_47# RESET_COUNTERn 0.01fF
C15216 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# SEL_CONV_TIME[0] 0.00fF
C15217 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C15218 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__inv_1_29/Y 0.00fF
C15219 DOUT[1] sky130_fd_sc_hd__dfrtn_1_23/a_639_47# 0.00fF
C15220 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C15221 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_543_47# 0.00fF
C15222 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_18/a_761_289# 0.00fF
C15223 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.00fF
C15224 sky130_fd_sc_hd__dfrtn_1_18/a_651_413# DOUT[2] 0.00fF
C15225 sky130_fd_sc_hd__o2111a_2_0/a_80_21# SEL_CONV_TIME[2] 0.00fF
C15226 sky130_fd_sc_hd__dfrtn_1_42/a_193_47# sky130_fd_sc_hd__inv_1_25/A 0.02fF
C15227 sky130_fd_sc_hd__dfrtn_1_32/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.02fF
C15228 sky130_fd_sc_hd__dfrtn_1_32/a_543_47# VDD 0.06fF
C15229 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# DOUT[11] 0.01fF
C15230 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C15231 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# -0.00fF
C15232 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C15233 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_448_47# -0.00fF
C15234 sky130_fd_sc_hd__dfrtn_1_36/a_761_289# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C15235 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__nand3b_1_0/Y 0.00fF
C15236 DOUT[16] sky130_fd_sc_hd__inv_1_52/Y -0.01fF
C15237 sky130_fd_sc_hd__dfrtn_1_36/a_193_47# sky130_fd_sc_hd__inv_1_52/Y 0.53fF
C15238 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# sky130_fd_sc_hd__inv_1_6/Y 0.01fF
C15239 sky130_fd_sc_hd__dfrtn_1_31/a_805_47# SEL_CONV_TIME[1] 0.00fF
C15240 DOUT[19] sky130_fd_sc_hd__inv_1_3/Y 0.05fF
C15241 sky130_fd_sc_hd__mux4_1_0/a_1290_413# RESET_COUNTERn 0.00fF
C15242 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_26/a_761_289# 0.00fF
C15243 sky130_fd_sc_hd__dfrtn_1_10/a_1217_47# RESET_COUNTERn 0.00fF
C15244 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_48/A 0.00fF
C15245 sky130_fd_sc_hd__dfrtn_1_21/a_1462_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C15246 sky130_fd_sc_hd__o211a_1_0/a_79_21# RESET_COUNTERn 0.01fF
C15247 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__dfrtn_1_28/a_27_47# 0.00fF
C15248 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_24/a_761_289# 0.01fF
C15249 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_19/a_1462_47# 0.00fF
C15250 sky130_fd_sc_hd__or3b_2_0/a_388_297# sky130_fd_sc_hd__dfrtn_1_31/a_448_47# 0.00fF
C15251 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_651_413# 0.00fF
C15252 sky130_fd_sc_hd__dfrtn_1_34/a_543_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C15253 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# 0.00fF
C15254 sky130_fd_sc_hd__dfrtn_1_28/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C15255 sky130_fd_sc_hd__dfrtn_1_17/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15256 sky130_fd_sc_hd__inv_1_39/A DOUT[15] 0.00fF
C15257 sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# VDD 0.00fF
C15258 sky130_fd_sc_hd__dfrtn_1_0/a_761_289# sky130_fd_sc_hd__nor3_1_0/a_193_297# 0.00fF
C15259 sky130_fd_sc_hd__dfrtn_1_0/a_543_47# sky130_fd_sc_hd__nor3_1_0/a_109_297# 0.00fF
C15260 sky130_fd_sc_hd__dfrtn_1_32/a_193_47# sky130_fd_sc_hd__dfrtn_1_32/a_448_47# -0.00fF
C15261 sky130_fd_sc_hd__dfrtn_1_32/a_27_47# sky130_fd_sc_hd__dfrtn_1_32/a_651_413# -0.00fF
C15262 HEADER_2/a_508_138# VDD 0.04fF
C15263 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# VDD 0.19fF
C15264 sky130_fd_sc_hd__dfrtn_1_22/a_651_413# sky130_fd_sc_hd__inv_1_37/A 0.01fF
C15265 sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C15266 DOUT[4] sky130_fd_sc_hd__dfrtn_1_30/a_193_47# 0.00fF
C15267 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# -0.00fF
C15268 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__dfrtn_1_30/a_543_47# -0.00fF
C15269 sky130_fd_sc_hd__nor3_1_0/A DOUT[17] 0.06fF
C15270 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C15271 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C15272 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C15273 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_448_47# 0.00fF
C15274 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__nor3_2_3/B 0.05fF
C15275 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# 0.00fF
C15276 sky130_fd_sc_hd__nor3_1_10/a_193_297# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C15277 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_1/A 0.01fF
C15278 sky130_fd_sc_hd__dfrtn_1_31/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15279 sky130_fd_sc_hd__dfrtn_1_31/a_639_47# VDD 0.00fF
C15280 sky130_fd_sc_hd__mux4_2_0/a_1064_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C15281 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__nor3_2_3/C 0.08fF
C15282 sky130_fd_sc_hd__mux4_2_0/a_1279_413# SEL_CONV_TIME[0] 0.00fF
C15283 sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C15284 sky130_fd_sc_hd__dfrtn_1_28/a_1283_21# sky130_fd_sc_hd__inv_1_42/A 0.00fF
C15285 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__mux4_1_0/X 0.01fF
C15286 sky130_fd_sc_hd__dfrtn_1_0/a_1462_47# RESET_COUNTERn 0.00fF
C15287 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C15288 sky130_fd_sc_hd__dfrtn_1_35/a_1270_413# RESET_COUNTERn 0.00fF
C15289 sky130_fd_sc_hd__nor3_1_4/a_109_297# DOUT[14] 0.00fF
C15290 sky130_fd_sc_hd__inv_1_32/A SEL_CONV_TIME[0] 0.01fF
C15291 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# sky130_fd_sc_hd__dfrtn_1_31/a_651_413# -0.00fF
C15292 sky130_fd_sc_hd__nor3_1_11/a_109_297# DOUT[6] 0.00fF
C15293 sky130_fd_sc_hd__nor3_1_11/a_193_297# DOUT[20] 0.00fF
C15294 sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C15295 sky130_fd_sc_hd__dfrtn_1_29/a_639_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C15296 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# 0.00fF
C15297 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_39/a_1462_47# 0.00fF
C15298 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_14/a_193_47# 0.00fF
C15299 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# RESET_COUNTERn 0.01fF
C15300 sky130_fd_sc_hd__dfrtn_1_4/a_651_413# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C15301 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# 0.00fF
C15302 sky130_fd_sc_hd__dfrtp_1_3/a_543_47# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C15303 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_543_47# 0.00fF
C15304 sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# sky130_fd_sc_hd__dfrtn_1_19/a_543_47# 0.00fF
C15305 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# sky130_fd_sc_hd__inv_1_31/A 0.00fF
C15306 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C15307 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__nor3_1_0/A 0.01fF
C15308 sky130_fd_sc_hd__inv_1_54/A sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# 0.00fF
C15309 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C15310 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_18/a_1462_47# 0.00fF
C15311 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_18/a_1270_413# 0.00fF
C15312 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_18/a_639_47# 0.00fF
C15313 sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C15314 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# 0.00fF
C15315 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C15316 sky130_fd_sc_hd__dfrtn_1_32/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15317 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__inv_1_7/A 0.61fF
C15318 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__dfrtn_1_29/a_761_289# 0.00fF
C15319 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C15320 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__dfrtn_1_29/a_543_47# 0.00fF
C15321 sky130_fd_sc_hd__dfrtn_1_10/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15322 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# CLK_REF 0.00fF
C15323 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C15324 sky130_fd_sc_hd__dfrtp_1_3/a_543_47# VDD 0.03fF
C15325 sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C15326 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_1/a_651_413# -0.00fF
C15327 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_1/a_448_47# -0.00fF
C15328 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# SEL_CONV_TIME[1] 0.00fF
C15329 sky130_fd_sc_hd__dfrtn_1_36/a_1462_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C15330 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_21/a_651_413# 0.00fF
C15331 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# sky130_fd_sc_hd__dfrtn_1_21/a_805_47# 0.00fF
C15332 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_1/A 0.00fF
C15333 sky130_fd_sc_hd__dfrtp_1_3/a_805_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C15334 sky130_fd_sc_hd__o311a_1_0/a_368_297# RESET_COUNTERn 0.00fF
C15335 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C15336 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C15337 sky130_fd_sc_hd__dfrtn_1_27/a_448_47# SEL_CONV_TIME[0] 0.00fF
C15338 sky130_fd_sc_hd__mux4_2_0/a_372_413# RESET_COUNTERn 0.00fF
C15339 sky130_fd_sc_hd__or2_2_0/a_121_297# RESET_COUNTERn 0.00fF
C15340 sky130_fd_sc_hd__or3_1_0/C sky130_fd_sc_hd__inv_1_48/Y 0.04fF
C15341 sky130_fd_sc_hd__inv_1_53/Y sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15342 sky130_fd_sc_hd__dfrtn_1_25/a_1462_47# sky130_fd_sc_hd__dfrtn_1_28/a_27_47# 0.00fF
C15343 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_36/a_651_413# 0.00fF
C15344 sky130_fd_sc_hd__dfrtn_1_24/a_1462_47# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C15345 sky130_fd_sc_hd__nor3_1_15/a_193_297# sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# 0.00fF
C15346 sky130_fd_sc_hd__nor3_1_8/a_193_297# DOUT[19] 0.00fF
C15347 sky130_fd_sc_hd__nor3_1_4/A RESET_COUNTERn 0.02fF
C15348 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_193_47# -0.17fF
C15349 sky130_fd_sc_hd__dfrtn_1_14/a_448_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C15350 sky130_fd_sc_hd__dfrtn_1_42/a_805_47# sky130_fd_sc_hd__nor3_2_3/A 0.00fF
C15351 sky130_fd_sc_hd__dfrtn_1_4/a_1270_413# DOUT[11] 0.00fF
C15352 sky130_fd_sc_hd__dfrtn_1_11/a_761_289# RESET_COUNTERn 0.01fF
C15353 sky130_fd_sc_hd__or2b_1_0/X sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C15354 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__o211a_1_1/X 0.01fF
C15355 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__dfrtn_1_33/a_1108_47# -0.00fF
C15356 sky130_fd_sc_hd__dfrtn_1_0/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15357 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15358 sky130_fd_sc_hd__dfrtn_1_14/a_639_47# DOUT[9] 0.00fF
C15359 sky130_fd_sc_hd__dfrtn_1_35/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15360 sky130_fd_sc_hd__nor3_1_20/a_109_297# RESET_COUNTERn 0.00fF
C15361 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# VDD 0.00fF
C15362 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C15363 sky130_fd_sc_hd__dfrtn_1_41/a_651_413# RESET_COUNTERn 0.01fF
C15364 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_34/a_1270_413# 0.00fF
C15365 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C15366 DOUT[4] sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# 0.00fF
C15367 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# VDD 0.10fF
C15368 sky130_fd_sc_hd__conb_1_0/LO DOUT[0] 0.00fF
C15369 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C15370 sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C15371 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C15372 sky130_fd_sc_hd__dfrtn_1_19/a_639_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C15373 sky130_fd_sc_hd__dfrtn_1_3/a_1270_413# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C15374 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__o211a_1_1/a_215_47# 0.00fF
C15375 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__o211a_1_1/a_297_297# 0.00fF
C15376 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__o211a_1_1/a_510_47# 0.00fF
C15377 sky130_fd_sc_hd__dfrtn_1_20/a_761_289# sky130_fd_sc_hd__dfrtn_1_18/a_193_47# 0.00fF
C15378 sky130_fd_sc_hd__dfrtn_1_20/a_543_47# sky130_fd_sc_hd__dfrtn_1_18/a_27_47# 0.01fF
C15379 sky130_fd_sc_hd__dfrtn_1_32/a_1270_413# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C15380 sky130_fd_sc_hd__dfrtp_1_2/a_448_47# sky130_fd_sc_hd__o211a_1_1/X 0.00fF
C15381 sky130_fd_sc_hd__inv_1_15/A RESET_COUNTERn 0.22fF
C15382 sky130_fd_sc_hd__dfrtn_1_23/a_761_289# sky130_fd_sc_hd__dfrtn_1_36/a_193_47# 0.00fF
C15383 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_543_47# 0.00fF
C15384 sky130_fd_sc_hd__dfrtn_1_23/a_543_47# sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C15385 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C15386 sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# DOUT[21] 0.00fF
C15387 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# RESET_COUNTERn 0.05fF
C15388 sky130_fd_sc_hd__dfrtn_1_38/a_193_47# sky130_fd_sc_hd__inv_1_53/A 0.03fF
C15389 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_21/a_543_47# 0.01fF
C15390 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# 0.00fF
C15391 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__or3_1_0/X 0.01fF
C15392 sky130_fd_sc_hd__dfrtn_1_35/a_193_47# sky130_fd_sc_hd__inv_1_38/A 0.01fF
C15393 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C15394 sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C15395 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__dfrtn_1_25/a_27_47# 0.00fF
C15396 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__dfrtn_1_25/a_448_47# 0.00fF
C15397 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__dfrtn_1_25/a_543_47# 0.00fF
C15398 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_32/a_543_47# 0.00fF
C15399 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C15400 sky130_fd_sc_hd__dfrtp_1_3/a_1217_47# sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# 0.00fF
C15401 sky130_fd_sc_hd__dfrtp_1_3/a_805_47# sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# 0.00fF
C15402 sky130_fd_sc_hd__inv_1_24/A DOUT[10] 0.00fF
C15403 sky130_fd_sc_hd__nor3_1_15/a_193_297# sky130_fd_sc_hd__dfrtn_1_32/a_193_47# 0.00fF
C15404 sky130_fd_sc_hd__o311a_1_0/a_81_21# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C15405 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__inv_1_6/Y 0.17fF
C15406 sky130_fd_sc_hd__dfrtn_1_12/a_1217_47# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C15407 sky130_fd_sc_hd__nor3_1_10/a_193_297# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C15408 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# sky130_fd_sc_hd__mux4_2_0/a_193_369# 0.00fF
C15409 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# sky130_fd_sc_hd__mux4_2_0/a_288_47# 0.00fF
C15410 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__mux4_2_0/a_600_345# 0.00fF
C15411 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# sky130_fd_sc_hd__mux4_2_0/a_788_316# 0.00fF
C15412 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C15413 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# sky130_fd_sc_hd__mux4_2_0/a_372_413# 0.00fF
C15414 sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C15415 sky130_fd_sc_hd__mux4_2_0/a_193_369# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15416 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C15417 sky130_fd_sc_hd__dfrtn_1_10/a_1283_21# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C15418 sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C15419 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# 0.00fF
C15420 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C15421 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C15422 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# 0.00fF
C15423 sky130_fd_sc_hd__o2111a_2_0/a_458_47# sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# 0.00fF
C15424 sky130_fd_sc_hd__a221oi_4_0/a_471_297# SEL_CONV_TIME[0] 0.01fF
C15425 sky130_fd_sc_hd__dfrtp_1_3/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15426 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# RESET_COUNTERn 0.03fF
C15427 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# 0.01fF
C15428 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# 0.00fF
C15429 sky130_fd_sc_hd__dfrtn_1_22/a_1108_47# VDD 0.07fF
C15430 sky130_fd_sc_hd__dfrtn_1_22/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15431 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C15432 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# RESET_COUNTERn 0.01fF
C15433 sky130_fd_sc_hd__dfrtn_1_20/a_543_47# sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# 0.00fF
C15434 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# -0.14fF
C15435 DOUT[1] sky130_fd_sc_hd__dfrtn_1_42/a_543_47# 0.00fF
C15436 sky130_fd_sc_hd__dfrtn_1_41/a_1270_413# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C15437 sky130_fd_sc_hd__dfrtn_1_28/a_651_413# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C15438 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__dfrtn_1_24/a_651_413# 0.00fF
C15439 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__inv_1_35/Y 0.02fF
C15440 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C15441 DOUT[4] sky130_fd_sc_hd__dfrtn_1_34/a_1270_413# 0.00fF
C15442 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# DOUT[2] 0.00fF
C15443 sky130_fd_sc_hd__nor3_1_13/a_193_297# outb 0.00fF
C15444 sky130_fd_sc_hd__or3b_2_0/a_176_21# SEL_CONV_TIME[0] 0.01fF
C15445 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__dfrtn_1_6/a_193_47# 0.00fF
C15446 sky130_fd_sc_hd__dfrtp_1_1/a_805_47# sky130_fd_sc_hd__dfrtp_1_1/D 0.00fF
C15447 sky130_fd_sc_hd__inv_1_33/A sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C15448 sky130_fd_sc_hd__dfrtn_1_23/a_448_47# sky130_fd_sc_hd__inv_1_40/A 0.00fF
C15449 sky130_fd_sc_hd__nand3b_1_0/a_316_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15450 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__dfrtp_1_1/a_193_47# 0.00fF
C15451 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/a_27_47# 0.00fF
C15452 sky130_fd_sc_hd__nand3b_1_1/a_232_47# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C15453 sky130_fd_sc_hd__inv_1_44/Y RESET_COUNTERn 0.12fF
C15454 sky130_fd_sc_hd__o311a_1_0/a_368_297# SEL_CONV_TIME[3] 0.00fF
C15455 sky130_fd_sc_hd__dfrtn_1_8/a_543_47# sky130_fd_sc_hd__inv_1_9/A 0.00fF
C15456 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_10/a_1270_413# 0.00fF
C15457 sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# DOUT[23] 0.00fF
C15458 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# DOUT[19] 0.00fF
C15459 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_48/A 0.03fF
C15460 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_543_47# 0.00fF
C15461 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_761_289# 0.00fF
C15462 sky130_fd_sc_hd__dfrtn_1_27/a_193_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C15463 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C15464 sky130_fd_sc_hd__dfrtn_1_8/a_1270_413# DOUT[12] 0.00fF
C15465 sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# sky130_fd_sc_hd__nor3_2_0/A 0.02fF
C15466 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C15467 sky130_fd_sc_hd__mux4_2_0/a_372_413# SEL_CONV_TIME[3] 0.00fF
C15468 sky130_fd_sc_hd__dfrtn_1_16/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.19fF
C15469 sky130_fd_sc_hd__dfrtn_1_16/a_543_47# VDD 0.06fF
C15470 sky130_fd_sc_hd__nor3_2_1/A sky130_fd_sc_hd__inv_1_26/A 0.00fF
C15471 SLC_0/a_264_22# sky130_fd_sc_hd__o211a_1_0/a_79_21# 0.00fF
C15472 sky130_fd_sc_hd__o211a_1_0/a_215_47# sky130_fd_sc_hd__inv_1_26/A 0.00fF
C15473 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15474 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C15475 sky130_fd_sc_hd__inv_1_14/A sky130_fd_sc_hd__nor3_1_5/a_193_297# 0.00fF
C15476 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__dfrtp_1_3/a_651_413# -0.00fF
C15477 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_448_47# -0.00fF
C15478 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# sky130_fd_sc_hd__inv_1_3/A 0.01fF
C15479 sky130_fd_sc_hd__a221oi_4_0/a_27_297# DOUT[21] 0.00fF
C15480 sky130_fd_sc_hd__inv_1_40/A DOUT[21] 0.06fF
C15481 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C15482 DOUT[9] sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C15483 CLK_REF sky130_fd_sc_hd__dfrtn_1_19/a_1270_413# 0.00fF
C15484 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15485 sky130_fd_sc_hd__dfrtn_1_20/a_1270_413# sky130_fd_sc_hd__dfrtn_1_18/a_448_47# 0.00fF
C15486 sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# sky130_fd_sc_hd__dfrtn_1_18/a_639_47# 0.00fF
C15487 sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# sky130_fd_sc_hd__dfrtn_1_18/a_805_47# 0.00fF
C15488 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C15489 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_20/a_193_47# 0.01fF
C15490 sky130_fd_sc_hd__dfrtn_1_18/a_651_413# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C15491 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__dfrtn_1_29/a_651_413# 0.00fF
C15492 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# SEL_CONV_TIME[0] 0.02fF
C15493 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C15494 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_40/a_761_289# -0.00fF
C15495 sky130_fd_sc_hd__dfrtp_1_0/a_1108_47# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C15496 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# sky130_fd_sc_hd__o211a_1_0/a_79_21# 0.00fF
C15497 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C15498 sky130_fd_sc_hd__dfrtn_1_23/a_1270_413# sky130_fd_sc_hd__dfrtn_1_36/a_448_47# 0.00fF
C15499 sky130_fd_sc_hd__dfrtn_1_23/a_1462_47# sky130_fd_sc_hd__dfrtn_1_36/a_761_289# 0.00fF
C15500 sky130_fd_sc_hd__dfrtn_1_23/a_1217_47# sky130_fd_sc_hd__dfrtn_1_36/a_543_47# 0.00fF
C15501 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# sky130_fd_sc_hd__dfrtn_1_36/a_805_47# 0.00fF
C15502 sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# sky130_fd_sc_hd__dfrtn_1_36/a_639_47# 0.00fF
C15503 sky130_fd_sc_hd__dfrtn_1_27/a_1217_47# RESET_COUNTERn 0.00fF
C15504 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# -0.00fF
C15505 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# -0.00fF
C15506 sky130_fd_sc_hd__dfrtn_1_26/a_761_289# sky130_fd_sc_hd__dfrtn_1_26/a_543_47# -0.00fF
C15507 sky130_fd_sc_hd__dfrtn_1_38/a_1462_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C15508 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15509 sky130_fd_sc_hd__dfrtn_1_35/a_1462_47# sky130_fd_sc_hd__inv_1_38/A 0.00fF
C15510 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C15511 sky130_fd_sc_hd__inv_1_26/A sky130_fd_sc_hd__or2_2_0/B 0.01fF
C15512 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C15513 sky130_fd_sc_hd__mux4_2_0/a_372_413# SEL_CONV_TIME[2] 0.00fF
C15514 sky130_fd_sc_hd__dfrtn_1_9/a_651_413# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C15515 sky130_fd_sc_hd__dfrtn_1_23/a_448_47# VDD 0.01fF
C15516 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15517 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_35/a_1108_47# 0.00fF
C15518 sky130_fd_sc_hd__dfrtn_1_30/a_639_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C15519 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__dfrtn_1_34/a_651_413# -0.00fF
C15520 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# sky130_fd_sc_hd__dfrtn_1_34/a_448_47# -0.00fF
C15521 DOUT[13] sky130_fd_sc_hd__dfrtn_1_30/a_651_413# 0.00fF
C15522 sky130_fd_sc_hd__dfrtn_1_38/a_805_47# DOUT[2] 0.00fF
C15523 sky130_fd_sc_hd__dfrtn_1_37/a_1462_47# sky130_fd_sc_hd__mux4_2_0/a_600_345# 0.00fF
C15524 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C15525 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# 0.00fF
C15526 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C15527 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C15528 sky130_fd_sc_hd__or3_1_0/C sky130_fd_sc_hd__nor3_2_3/B 0.24fF
C15529 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15530 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# VDD 0.03fF
C15531 sky130_fd_sc_hd__mux4_2_0/a_1281_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15532 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__inv_1_15/A 0.00fF
C15533 sky130_fd_sc_hd__dfrtn_1_36/a_543_47# RESET_COUNTERn 0.02fF
C15534 sky130_fd_sc_hd__dfrtn_1_36/a_1270_413# DOUT[21] 0.00fF
C15535 sky130_fd_sc_hd__dfrtn_1_37/a_1270_413# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C15536 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C15537 CLK_REF sky130_fd_sc_hd__inv_1_34/A 0.06fF
C15538 DOUT[4] sky130_fd_sc_hd__dfrtn_1_28/a_193_47# 0.00fF
C15539 sky130_fd_sc_hd__dfrtp_1_0/a_1108_47# sky130_fd_sc_hd__or2_2_0/B 0.01fF
C15540 sky130_fd_sc_hd__dfrtn_1_9/a_805_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C15541 sky130_fd_sc_hd__o311a_1_0/a_81_21# sky130_fd_sc_hd__nand2_1_1/Y 0.05fF
C15542 sky130_fd_sc_hd__or2b_1_0/X sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C15543 sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C15544 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# VDD 0.00fF
C15545 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15546 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C15547 sky130_fd_sc_hd__dfrtn_1_11/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15548 VDD DOUT[21] 2.12fF
C15549 sky130_fd_sc_hd__nor3_1_12/a_193_297# sky130_fd_sc_hd__dfrtn_1_8/a_651_413# 0.00fF
C15550 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C15551 sky130_fd_sc_hd__nand2_1_1/a_113_47# SEL_CONV_TIME[3] 0.00fF
C15552 sky130_fd_sc_hd__dfrtn_1_18/a_27_47# sky130_fd_sc_hd__inv_1_35/A 0.00fF
C15553 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__inv_1_47/Y 0.00fF
C15554 sky130_fd_sc_hd__dfrtn_1_21/a_651_413# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C15555 sky130_fd_sc_hd__dfrtn_1_18/a_805_47# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C15556 sky130_fd_sc_hd__o2111a_2_0/a_458_47# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C15557 sky130_fd_sc_hd__nor3_1_7/a_109_297# RESET_COUNTERn 0.00fF
C15558 sky130_fd_sc_hd__dfrtn_1_27/a_543_47# DOUT[23] 0.00fF
C15559 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# 0.00fF
C15560 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# 0.00fF
C15561 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# 0.00fF
C15562 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__or3_1_0/C 0.01fF
C15563 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__mux4_2_0/a_1281_47# 0.00fF
C15564 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# DOUT[0] 0.00fF
C15565 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C15566 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# 0.01fF
C15567 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_543_47# 0.01fF
C15568 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.00fF
C15569 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# sky130_fd_sc_hd__nor3_1_4/A 0.01fF
C15570 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__dfrtn_1_13/a_543_47# 0.00fF
C15571 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C15572 sky130_fd_sc_hd__dfrtn_1_26/a_448_47# sky130_fd_sc_hd__dfrtn_1_38/a_1270_413# 0.00fF
C15573 sky130_fd_sc_hd__dfrtn_1_42/a_761_289# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C15574 sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C15575 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C15576 sky130_fd_sc_hd__dfrtn_1_16/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15577 sky130_fd_sc_hd__dfrtn_1_27/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15578 sky130_fd_sc_hd__dfrtn_1_8/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15579 sky130_fd_sc_hd__dfrtn_1_8/a_805_47# VDD 0.00fF
C15580 VDD sky130_fd_sc_hd__o311a_1_0/A3 0.22fF
C15581 sky130_fd_sc_hd__nand2_1_1/a_113_47# SEL_CONV_TIME[2] 0.00fF
C15582 sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# sky130_fd_sc_hd__inv_1_49/A 0.02fF
C15583 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C15584 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_639_47# -0.00fF
C15585 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__inv_1_7/A 0.01fF
C15586 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C15587 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C15588 sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# DOUT[21] 0.00fF
C15589 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C15590 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__dfrtn_1_34/a_193_47# 0.00fF
C15591 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__dfrtn_1_34/a_761_289# 0.00fF
C15592 sky130_fd_sc_hd__inv_1_44/Y SEL_CONV_TIME[3] 0.02fF
C15593 sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# sky130_fd_sc_hd__inv_1_35/A 0.01fF
C15594 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_20/a_1462_47# 0.00fF
C15595 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# CLK_REF 0.02fF
C15596 DOUT[4] sky130_fd_sc_hd__dfrtn_1_10/a_1283_21# 0.00fF
C15597 sky130_fd_sc_hd__dfrtn_1_31/a_1217_47# SEL_CONV_TIME[0] 0.00fF
C15598 sky130_fd_sc_hd__o311a_1_0/a_266_297# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C15599 DOUT[16] sky130_fd_sc_hd__nor3_2_3/B 0.08fF
C15600 sky130_fd_sc_hd__dfrtn_1_36/a_193_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15601 sky130_fd_sc_hd__inv_1_22/Y sky130_fd_sc_hd__inv_1_23/A 0.03fF
C15602 HEADER_0/a_508_138# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C15603 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15604 sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C15605 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# sky130_fd_sc_hd__inv_1_44/A 0.01fF
C15606 sky130_fd_sc_hd__nor3_1_4/A DOUT[10] 0.01fF
C15607 sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C15608 sky130_fd_sc_hd__dfrtn_1_25/a_448_47# sky130_fd_sc_hd__or3_1_0/C 0.01fF
C15609 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__nor3_2_0/A 0.02fF
C15610 sky130_fd_sc_hd__dfrtn_1_12/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15611 sky130_fd_sc_hd__nor3_2_0/a_281_297# VDD 0.04fF
C15612 sky130_fd_sc_hd__dfrtn_1_39/a_761_289# sky130_fd_sc_hd__inv_1_32/A 0.01fF
C15613 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__mux4_2_0/a_193_47# 0.00fF
C15614 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# 0.00fF
C15615 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_3/a_805_47# 0.00fF
C15616 sky130_fd_sc_hd__dfrtn_1_7/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15617 sky130_fd_sc_hd__dfrtn_1_17/a_651_413# RESET_COUNTERn 0.00fF
C15618 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# DOUT[14] 0.00fF
C15619 sky130_fd_sc_hd__dfrtn_1_41/a_448_47# sky130_fd_sc_hd__inv_1_54/A 0.00fF
C15620 sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C15621 sky130_fd_sc_hd__or2_2_0/A sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C15622 DOUT[6] DOUT[14] 0.04fF
C15623 sky130_fd_sc_hd__dfrtn_1_9/a_639_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C15624 DOUT[4] sky130_fd_sc_hd__dfrtn_1_28/a_1462_47# 0.00fF
C15625 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__inv_1_7/A 0.01fF
C15626 sky130_fd_sc_hd__nor3_1_1/a_193_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15627 sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# sky130_fd_sc_hd__inv_1_0/Y 0.01fF
C15628 DOUT[4] sky130_fd_sc_hd__dfrtn_1_35/a_193_47# 0.01fF
C15629 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# sky130_fd_sc_hd__inv_1_11/Y 0.01fF
C15630 sky130_fd_sc_hd__inv_1_27/Y sky130_fd_sc_hd__inv_1_53/A 0.09fF
C15631 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_651_413# 0.00fF
C15632 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# 0.00fF
C15633 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_2/a_761_289# 0.00fF
C15634 sky130_fd_sc_hd__dfrtn_1_31/a_1108_47# RESET_COUNTERn -0.00fF
C15635 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C15636 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C15637 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C15638 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_12/a_27_47# 0.02fF
C15639 sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C15640 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# SEL_CONV_TIME[1] 0.01fF
C15641 sky130_fd_sc_hd__nor3_1_13/a_193_297# sky130_fd_sc_hd__dfrtn_1_10/a_448_47# 0.00fF
C15642 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C15643 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.00fF
C15644 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C15645 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C15646 sky130_fd_sc_hd__dfrtn_1_25/a_651_413# sky130_fd_sc_hd__dfrtn_1_27/a_1270_413# 0.00fF
C15647 sky130_fd_sc_hd__dfrtn_1_25/a_805_47# sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# 0.00fF
C15648 sky130_fd_sc_hd__dfrtn_1_25/a_1217_47# sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# 0.00fF
C15649 sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# DOUT[2] 0.01fF
C15650 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__dfrtn_1_23/a_193_47# 0.00fF
C15651 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# sky130_fd_sc_hd__dfrtn_1_23/a_27_47# 0.00fF
C15652 sky130_fd_sc_hd__dfrtn_1_31/a_543_47# DONE 0.00fF
C15653 sky130_fd_sc_hd__mux4_2_0/a_193_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C15654 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_21/a_639_47# 0.00fF
C15655 sky130_fd_sc_hd__dfrtn_1_9/a_761_289# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C15656 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__inv_1_27/Y 0.04fF
C15657 sky130_fd_sc_hd__or3b_2_0/a_472_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15658 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C15659 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C15660 VDD sky130_fd_sc_hd__dfrtp_1_1/D 0.13fF
C15661 sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C15662 sky130_fd_sc_hd__dfrtn_1_23/a_1217_47# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C15663 sky130_fd_sc_hd__dfrtn_1_32/a_805_47# RESET_COUNTERn 0.00fF
C15664 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# SEL_CONV_TIME[0] 0.00fF
C15665 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__dfrtn_1_33/a_193_47# 0.00fF
C15666 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__dfrtn_1_33/a_761_289# 0.00fF
C15667 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__dfrtn_1_33/a_543_47# 0.00fF
C15668 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_33/a_448_47# 0.00fF
C15669 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_33/a_27_47# 0.00fF
C15670 sky130_fd_sc_hd__o311a_1_0/a_368_297# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C15671 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# sky130_fd_sc_hd__dfrtn_1_14/a_448_47# -0.00fF
C15672 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# sky130_fd_sc_hd__dfrtn_1_14/a_651_413# -0.00fF
C15673 sky130_fd_sc_hd__dfrtn_1_8/a_639_47# sky130_fd_sc_hd__inv_1_9/Y 0.00fF
C15674 sky130_fd_sc_hd__dfrtn_1_28/a_1270_413# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C15675 sky130_fd_sc_hd__or3_1_0/a_111_297# sky130_fd_sc_hd__a221oi_4_0/a_1241_47# 0.00fF
C15676 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C15677 sky130_fd_sc_hd__dfrtn_1_10/a_1283_21# outb 0.00fF
C15678 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# sky130_fd_sc_hd__dfrtn_1_22/a_805_47# -0.00fF
C15679 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# sky130_fd_sc_hd__dfrtn_1_22/a_1217_47# -0.00fF
C15680 sky130_fd_sc_hd__dfrtn_1_36/a_1462_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15681 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__o211a_1_1/X 0.00fF
C15682 sky130_fd_sc_hd__inv_1_25/A sky130_fd_sc_hd__nor3_2_3/A 0.14fF
C15683 sky130_fd_sc_hd__or2b_1_0/a_301_297# RESET_COUNTERn 0.00fF
C15684 sky130_fd_sc_hd__dfrtn_1_37/a_639_47# VDD 0.00fF
C15685 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C15686 sky130_fd_sc_hd__inv_1_52/Y RESET_COUNTERn 0.24fF
C15687 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_17/a_805_47# 0.00fF
C15688 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__inv_1_46/Y 0.00fF
C15689 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15690 sky130_fd_sc_hd__dfrtn_1_3/a_1270_413# VDD 0.00fF
C15691 sky130_fd_sc_hd__dfrtn_1_14/a_448_47# sky130_fd_sc_hd__inv_1_1/A 0.01fF
C15692 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# 0.00fF
C15693 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# 0.00fF
C15694 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__dfrtp_1_2/a_193_47# 0.00fF
C15695 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_2/a_543_47# 0.00fF
C15696 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__dfrtp_1_2/a_761_289# 0.00fF
C15697 sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C15698 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C15699 sky130_fd_sc_hd__inv_1_10/A DOUT[21] 0.55fF
C15700 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C15701 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C15702 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C15703 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# 0.01fF
C15704 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C15705 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_448_47# 0.00fF
C15706 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_5/A 0.00fF
C15707 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C15708 DOUT[2] sky130_fd_sc_hd__inv_1_53/Y 0.03fF
C15709 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# RESET_COUNTERn 0.00fF
C15710 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# VDD 0.18fF
C15711 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C15712 sky130_fd_sc_hd__dfrtn_1_19/a_805_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C15713 DOUT[4] sky130_fd_sc_hd__dfrtn_1_35/a_1462_47# 0.00fF
C15714 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# 0.00fF
C15715 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# DOUT[21] 0.00fF
C15716 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# RESET_COUNTERn 0.29fF
C15717 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_31/a_1270_413# 0.00fF
C15718 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C15719 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__dfrtn_1_23/a_761_289# -0.00fF
C15720 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__inv_1_37/A 0.02fF
C15721 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C15722 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# VDD 0.06fF
C15723 sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C15724 sky130_fd_sc_hd__dfrtn_1_4/a_761_289# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C15725 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15726 sky130_fd_sc_hd__dfrtn_1_38/a_761_289# sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C15727 sky130_fd_sc_hd__dfrtn_1_14/a_761_289# DOUT[11] 0.00fF
C15728 sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# VDD 0.10fF
C15729 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C15730 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# 0.00fF
C15731 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__nor3_2_3/B 0.03fF
C15732 sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# 0.00fF
C15733 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__dfrtn_1_26/a_651_413# 0.00fF
C15734 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_26/a_27_47# 0.00fF
C15735 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__dfrtn_1_26/a_639_47# 0.00fF
C15736 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# DOUT[3] 0.00fF
C15737 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_29/a_761_289# 0.00fF
C15738 sky130_fd_sc_hd__dfrtn_1_32/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15739 sky130_fd_sc_hd__dfrtn_1_25/a_1217_47# SEL_CONV_TIME[1] 0.00fF
C15740 sky130_fd_sc_hd__dfrtn_1_21/a_651_413# VDD 0.01fF
C15741 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C15742 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_8/a_805_47# 0.00fF
C15743 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# 0.00fF
C15744 sky130_fd_sc_hd__dfrtn_1_19/a_651_413# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C15745 sky130_fd_sc_hd__o211a_1_1/a_215_47# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C15746 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# sky130_fd_sc_hd__dfrtn_1_16/a_651_413# -0.00fF
C15747 sky130_fd_sc_hd__dfrtn_1_16/a_193_47# sky130_fd_sc_hd__dfrtn_1_16/a_448_47# -0.00fF
C15748 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C15749 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# DOUT[3] 0.00fF
C15750 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# DOUT[2] 0.00fF
C15751 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# sky130_fd_sc_hd__o311a_1_0/A3 0.02fF
C15752 sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# sky130_fd_sc_hd__inv_1_27/Y 0.00fF
C15753 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_27_47# 0.01fF
C15754 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C15755 sky130_fd_sc_hd__nor3_1_20/a_109_297# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C15756 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__nor3_1_4/a_109_297# 0.00fF
C15757 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_3/a_761_289# 0.00fF
C15758 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_0/a_543_47# 0.02fF
C15759 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15760 sky130_fd_sc_hd__nor3_2_2/a_281_297# sky130_fd_sc_hd__dfrtn_1_16/a_1108_47# 0.00fF
C15761 sky130_fd_sc_hd__mux4_2_0/a_372_413# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C15762 sky130_fd_sc_hd__dfrtn_1_28/a_193_47# sky130_fd_sc_hd__dfrtn_1_28/a_543_47# -0.00fF
C15763 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C15764 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C15765 sky130_fd_sc_hd__dfrtp_1_0/a_761_289# VDD 0.05fF
C15766 sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# sky130_fd_sc_hd__or2_2_0/X 0.00fF
C15767 sky130_fd_sc_hd__dfrtp_1_3/a_805_47# RESET_COUNTERn 0.00fF
C15768 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# -0.00fF
C15769 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1_6/a_448_47# -0.00fF
C15770 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# sky130_fd_sc_hd__o211a_1_1/a_215_47# 0.00fF
C15771 sky130_fd_sc_hd__dfrtp_1_1/a_639_47# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.00fF
C15772 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C15773 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C15774 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# RESET_COUNTERn 0.00fF
C15775 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_761_289# 0.01fF
C15776 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C15777 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C15778 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C15779 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.01fF
C15780 sky130_fd_sc_hd__dfrtn_1_39/a_543_47# VDD 0.10fF
C15781 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15782 sky130_fd_sc_hd__dfrtn_1_25/a_805_47# VDD 0.00fF
C15783 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__nor3_2_0/a_281_297# 0.00fF
C15784 sky130_fd_sc_hd__dfrtn_1_41/a_651_413# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C15785 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__dfrtn_1_3/a_27_47# 0.00fF
C15786 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_3/a_448_47# 0.00fF
C15787 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# sky130_fd_sc_hd__dfrtn_1_3/a_651_413# 0.00fF
C15788 sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# sky130_fd_sc_hd__dfrtn_1_3/a_193_47# 0.00fF
C15789 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# 0.00fF
C15790 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# 0.00fF
C15791 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_639_47# 0.00fF
C15792 sky130_fd_sc_hd__or3_1_0/X sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C15793 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C15794 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# sky130_fd_sc_hd__nor3_1_5/a_193_297# 0.00fF
C15795 sky130_fd_sc_hd__o221ai_1_0/a_493_297# SEL_CONV_TIME[1] 0.00fF
C15796 sky130_fd_sc_hd__dfrtn_1_18/a_543_47# VDD 0.06fF
C15797 sky130_fd_sc_hd__dfrtn_1_20/a_639_47# sky130_fd_sc_hd__inv_1_35/Y 0.00fF
C15798 DOUT[9] VDD 2.66fF
C15799 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__inv_1_5/Y 0.01fF
C15800 sky130_fd_sc_hd__inv_1_45/Y DOUT[2] 0.00fF
C15801 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# DOUT[2] 0.00fF
C15802 sky130_fd_sc_hd__dfrtn_1_24/a_805_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C15803 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C15804 sky130_fd_sc_hd__dfrtn_1_24/a_1270_413# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C15805 sky130_fd_sc_hd__dfrtn_1_42/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15806 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__nor3_2_1/a_27_297# 0.00fF
C15807 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__nor3_2_1/a_281_297# 0.00fF
C15808 sky130_fd_sc_hd__dfrtn_1_42/a_1217_47# VDD 0.00fF
C15809 sky130_fd_sc_hd__inv_1_11/A sky130_fd_sc_hd__inv_1_5/A 0.00fF
C15810 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__nor3_2_3/B 0.14fF
C15811 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__inv_1_29/Y 0.00fF
C15812 sky130_fd_sc_hd__dfrtn_1_8/a_27_47# DOUT[21] 0.01fF
C15813 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# DOUT[14] 0.01fF
C15814 sky130_fd_sc_hd__dfrtn_1_4/a_448_47# DOUT[14] 0.00fF
C15815 sky130_fd_sc_hd__nor3_1_5/a_193_297# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C15816 VDD sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.07fF
C15817 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# 0.00fF
C15818 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C15819 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C15820 sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# RESET_COUNTERn 0.00fF
C15821 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C15822 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_25/a_448_47# 0.00fF
C15823 sky130_fd_sc_hd__dfrtn_1_38/a_761_289# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C15824 sky130_fd_sc_hd__dfrtn_1_10/a_805_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C15825 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# 0.00fF
C15826 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_38/a_651_413# 0.00fF
C15827 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# sky130_fd_sc_hd__dfrtn_1_38/a_761_289# 0.00fF
C15828 sky130_fd_sc_hd__dfrtn_1_41/a_651_413# sky130_fd_sc_hd__dfrtn_1_38/a_27_47# 0.00fF
C15829 sky130_fd_sc_hd__dfrtn_1_41/a_448_47# sky130_fd_sc_hd__dfrtn_1_38/a_193_47# 0.00fF
C15830 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# sky130_fd_sc_hd__dfrtn_1_38/a_448_47# 0.00fF
C15831 sky130_fd_sc_hd__dfrtp_1_3/a_761_289# DOUT[23] 0.00fF
C15832 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# VDD 0.00fF
C15833 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15834 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__inv_1_43/Y 0.08fF
C15835 sky130_fd_sc_hd__nor3_1_3/a_193_297# RESET_COUNTERn 0.00fF
C15836 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# 0.00fF
C15837 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__dfrtn_1_1/a_27_47# 0.00fF
C15838 sky130_fd_sc_hd__o311a_1_0/a_266_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C15839 sky130_fd_sc_hd__o221ai_1_0/a_295_297# VDD 0.00fF
C15840 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C15841 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C15842 sky130_fd_sc_hd__inv_1_22/Y DOUT[10] 0.01fF
C15843 sky130_fd_sc_hd__inv_1_3/A sky130_fd_sc_hd__inv_1_2/Y 0.01fF
C15844 sky130_fd_sc_hd__nor3_1_4/A sky130_fd_sc_hd__inv_1_4/Y 0.09fF
C15845 sky130_fd_sc_hd__nor3_1_14/a_193_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15846 sky130_fd_sc_hd__dfrtn_1_19/a_448_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C15847 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__inv_1_41/Y 0.01fF
C15848 sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# SEL_CONV_TIME[1] 0.01fF
C15849 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# SEL_CONV_TIME[3] 0.00fF
C15850 sky130_fd_sc_hd__dfrtp_1_3/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15851 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# sky130_fd_sc_hd__dfrtn_1_7/a_543_47# -0.00fF
C15852 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# -0.00fF
C15853 sky130_fd_sc_hd__inv_1_49/Y SEL_CONV_TIME[1] 0.02fF
C15854 sky130_fd_sc_hd__dfrtn_1_16/a_651_413# DOUT[15] 0.01fF
C15855 sky130_fd_sc_hd__dfrtn_1_33/a_448_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C15856 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C15857 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C15858 DOUT[11] sky130_fd_sc_hd__inv_1_7/A 0.01fF
C15859 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C15860 sky130_fd_sc_hd__dfrtn_1_23/a_651_413# DOUT[21] 0.00fF
C15861 sky130_fd_sc_hd__dfrtn_1_23/a_761_289# RESET_COUNTERn 0.01fF
C15862 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C15863 sky130_fd_sc_hd__dfrtn_1_41/a_1270_413# sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.00fF
C15864 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# 0.00fF
C15865 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# sky130_fd_sc_hd__dfrtn_1_7/a_805_47# 0.00fF
C15866 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# sky130_fd_sc_hd__dfrtn_1_7/a_761_289# 0.00fF
C15867 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# sky130_fd_sc_hd__dfrtn_1_7/a_448_47# 0.00fF
C15868 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# sky130_fd_sc_hd__dfrtn_1_7/a_543_47# 0.00fF
C15869 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__dfrtn_1_7/a_1217_47# 0.00fF
C15870 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# sky130_fd_sc_hd__dfrtn_1_7/a_193_47# 0.00fF
C15871 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# sky130_fd_sc_hd__dfrtn_1_7/a_639_47# 0.00fF
C15872 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# sky130_fd_sc_hd__dfrtn_1_7/a_27_47# 0.00fF
C15873 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# 0.00fF
C15874 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C15875 DOUT[4] sky130_fd_sc_hd__dfrtn_1_12/a_651_413# 0.00fF
C15876 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# sky130_fd_sc_hd__inv_1_11/A 0.00fF
C15877 sky130_fd_sc_hd__dfrtn_1_12/a_651_413# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C15878 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# DOUT[20] 0.01fF
C15879 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# DOUT[7] 0.02fF
C15880 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# DOUT[6] 0.01fF
C15881 sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C15882 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/X 0.01fF
C15883 sky130_fd_sc_hd__dfrtp_1_0/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15884 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_0/a_193_47# -0.32fF
C15885 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# DOUT[6] 0.00fF
C15886 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# RESET_COUNTERn 0.01fF
C15887 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# DOUT[7] 0.00fF
C15888 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# DOUT[8] 0.00fF
C15889 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# DOUT[20] 0.00fF
C15890 DOUT[22] DOUT[18] 0.02fF
C15891 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__inv_1_43/A 0.03fF
C15892 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_2/Y 0.29fF
C15893 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C15894 sky130_fd_sc_hd__inv_1_53/A sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C15895 sky130_fd_sc_hd__dfrtn_1_22/a_1462_47# RESET_COUNTERn 0.00fF
C15896 sky130_fd_sc_hd__inv_1_21/Y sky130_fd_sc_hd__inv_1_19/A 0.00fF
C15897 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C15898 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.00fF
C15899 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C15900 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# 0.00fF
C15901 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# 0.00fF
C15902 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# SEL_CONV_TIME[2] 0.00fF
C15903 CLK_REF sky130_fd_sc_hd__dfrtn_1_20/a_639_47# 0.00fF
C15904 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_32/a_651_413# 0.00fF
C15905 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C15906 sky130_fd_sc_hd__o2111a_2_0/a_566_47# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C15907 sky130_fd_sc_hd__dfrtn_1_31/a_448_47# sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C15908 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# sky130_fd_sc_hd__inv_1_42/Y 0.01fF
C15909 sky130_fd_sc_hd__dfrtn_1_26/a_761_289# sky130_fd_sc_hd__dfrtn_1_27/a_27_47# 0.00fF
C15910 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.00fF
C15911 sky130_fd_sc_hd__inv_1_48/Y RESET_COUNTERn 0.03fF
C15912 sky130_fd_sc_hd__dfrtn_1_30/a_639_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C15913 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15914 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# VDD 0.06fF
C15915 sky130_fd_sc_hd__o2111a_2_0/a_80_21# sky130_fd_sc_hd__o311a_1_0/a_266_297# 0.00fF
C15916 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.00fF
C15917 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_10/a_805_47# -0.00fF
C15918 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__inv_1_32/A 0.01fF
C15919 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# outb 0.00fF
C15920 sky130_fd_sc_hd__nor3_1_19/Y sky130_fd_sc_hd__inv_1_33/A 0.00fF
C15921 sky130_fd_sc_hd__dfrtn_1_29/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15922 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# SEL_CONV_TIME[0] 0.00fF
C15923 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__dfrtn_1_3/a_193_47# 0.00fF
C15924 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__dfrtn_1_3/a_27_47# 0.00fF
C15925 sky130_fd_sc_hd__dfrtn_1_9/a_761_289# DOUT[14] 0.00fF
C15926 sky130_fd_sc_hd__nor3_1_19/a_193_297# sky130_fd_sc_hd__mux4_2_0/a_27_47# 0.00fF
C15927 sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# sky130_fd_sc_hd__dfrtn_1_19/a_448_47# 0.00fF
C15928 sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# sky130_fd_sc_hd__dfrtn_1_19/a_651_413# 0.00fF
C15929 sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C15930 sky130_fd_sc_hd__dfrtn_1_26/a_448_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C15931 sky130_fd_sc_hd__dfrtn_1_16/a_805_47# RESET_COUNTERn 0.00fF
C15932 sky130_fd_sc_hd__dfrtn_1_8/a_448_47# RESET_COUNTERn 0.00fF
C15933 sky130_fd_sc_hd__dfrtn_1_8/a_1217_47# DOUT[21] 0.00fF
C15934 sky130_fd_sc_hd__or3b_2_0/B SEL_CONV_TIME[0] 0.03fF
C15935 DOUT[4] SEL_CONV_TIME[1] 0.11fF
C15936 sky130_fd_sc_hd__dfrtp_1_0/a_761_289# sky130_fd_sc_hd__o211a_1_0/X 0.00fF
C15937 sky130_fd_sc_hd__dfrtn_1_9/a_639_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15938 VDD sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# 0.00fF
C15939 sky130_fd_sc_hd__dfrtn_1_30/a_543_47# SEL_CONV_TIME[1] 0.01fF
C15940 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# sky130_fd_sc_hd__dfrtn_1_20/a_1217_47# -0.00fF
C15941 sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C15942 sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# sky130_fd_sc_hd__inv_1_36/Y 0.00fF
C15943 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15944 sky130_fd_sc_hd__dfrtn_1_19/a_805_47# VDD 0.00fF
C15945 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# 0.00fF
C15946 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_30/a_27_47# 0.00fF
C15947 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_30/a_193_47# 0.00fF
C15948 sky130_fd_sc_hd__nor3_1_8/a_109_297# VDD 0.00fF
C15949 sky130_fd_sc_hd__nor3_1_0/a_193_297# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C15950 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C15951 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__dfrtn_1_1/a_448_47# 0.00fF
C15952 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__dfrtn_1_1/a_805_47# 0.00fF
C15953 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C15954 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__dfrtn_1_18/a_805_47# 0.00fF
C15955 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C15956 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__inv_1_48/A 0.01fF
C15957 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C15958 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C15959 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_27/a_651_413# 0.00fF
C15960 DOUT[4] sky130_fd_sc_hd__dfrtn_1_36/a_651_413# 0.00fF
C15961 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15962 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# 0.00fF
C15963 sky130_fd_sc_hd__dfrtn_1_22/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15964 sky130_fd_sc_hd__nor3_1_3/a_193_297# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C15965 sky130_fd_sc_hd__dfrtn_1_7/a_1217_47# DOUT[7] 0.00fF
C15966 sky130_fd_sc_hd__dfrtn_1_7/a_639_47# RESET_COUNTERn 0.00fF
C15967 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15968 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# DOUT[3] 0.00fF
C15969 sky130_fd_sc_hd__dfrtn_1_30/a_761_289# VDD 0.06fF
C15970 sky130_fd_sc_hd__inv_1_54/Y sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C15971 sky130_fd_sc_hd__inv_1_47/Y SEL_CONV_TIME[1] 0.02fF
C15972 sky130_fd_sc_hd__dfrtn_1_30/a_448_47# sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.00fF
C15973 sky130_fd_sc_hd__dfrtn_1_16/a_761_289# DOUT[23] 0.00fF
C15974 sky130_fd_sc_hd__dfrtn_1_14/a_448_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C15975 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# sky130_fd_sc_hd__dfrtn_1_31/a_27_47# 0.00fF
C15976 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# sky130_fd_sc_hd__dfrtn_1_31/a_193_47# 0.00fF
C15977 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# DOUT[14] 0.02fF
C15978 sky130_fd_sc_hd__dfrtn_1_14/a_543_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C15979 sky130_fd_sc_hd__dfrtn_1_35/a_193_47# sky130_fd_sc_hd__dfrtn_1_35/a_543_47# -0.00fF
C15980 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# sky130_fd_sc_hd__dfrtn_1_35/a_1283_21# -0.00fF
C15981 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_2/A 0.01fF
C15982 sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# CLK_REF 0.00fF
C15983 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C15984 sky130_fd_sc_hd__nor3_1_3/a_109_297# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C15985 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__inv_1_39/Y 0.01fF
C15986 sky130_fd_sc_hd__nor3_2_0/A sky130_fd_sc_hd__inv_1_5/A 0.00fF
C15987 sky130_fd_sc_hd__dfrtn_1_14/a_448_47# DOUT[17] 0.00fF
C15988 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_1290_413# -0.00fF
C15989 sky130_fd_sc_hd__dfrtn_1_27/a_1217_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C15990 sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.00fF
C15991 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# sky130_fd_sc_hd__dfrtn_1_27/a_639_47# 0.00fF
C15992 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C15993 sky130_fd_sc_hd__nor3_2_2/a_281_297# DOUT[23] 0.00fF
C15994 sky130_fd_sc_hd__dfrtn_1_24/a_1462_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15995 sky130_fd_sc_hd__dfrtn_1_16/a_1270_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C15996 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C15997 sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C15998 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# SEL_CONV_TIME[0] 0.00fF
C15999 lc_out RESET_COUNTERn 0.02fF
C16000 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# VDD 0.00fF
C16001 sky130_fd_sc_hd__dfrtn_1_8/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C16002 sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C16003 sky130_fd_sc_hd__inv_1_36/A sky130_fd_sc_hd__inv_1_9/A 0.00fF
C16004 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C16005 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_11/a_27_47# 0.00fF
C16006 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_193_47# 0.00fF
C16007 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C16008 DONE RESET_COUNTERn 0.01fF
C16009 sky130_fd_sc_hd__nor3_1_17/a_193_297# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C16010 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# 0.01fF
C16011 sky130_fd_sc_hd__o2111a_2_0/a_674_297# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C16012 DOUT[4] sky130_fd_sc_hd__dfrtn_1_32/a_543_47# 0.00fF
C16013 sky130_fd_sc_hd__dfrtn_1_12/a_761_289# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C16014 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__dfrtn_1_40/a_27_47# 0.00fF
C16015 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__dfrtn_1_40/a_193_47# 0.00fF
C16016 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# 0.00fF
C16017 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_17/a_193_47# 0.00fF
C16018 sky130_fd_sc_hd__dfrtp_1_2/a_448_47# sky130_fd_sc_hd__dfrtn_1_17/a_27_47# 0.00fF
C16019 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_448_47# 0.00fF
C16020 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__dfrtn_1_17/a_543_47# 0.00fF
C16021 sky130_fd_sc_hd__dfrtn_1_12/a_761_289# sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# 0.00fF
C16022 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# 0.00fF
C16023 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# sky130_fd_sc_hd__dfrtn_1_14/a_27_47# 0.00fF
C16024 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_14/a_27_47# 0.02fF
C16025 sky130_fd_sc_hd__nor3_2_2/a_27_297# sky130_fd_sc_hd__dfrtn_1_42/a_543_47# 0.00fF
C16026 sky130_fd_sc_hd__nor3_1_19/a_109_297# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C16027 sky130_fd_sc_hd__dfrtn_1_20/a_651_413# sky130_fd_sc_hd__dfrtn_1_21/a_27_47# 0.00fF
C16028 sky130_fd_sc_hd__dfrtn_1_23/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C16029 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# sky130_fd_sc_hd__inv_1_6/A 0.01fF
C16030 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# DOUT[14] 0.01fF
C16031 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# sky130_fd_sc_hd__inv_1_30/Y 0.00fF
C16032 sky130_fd_sc_hd__nor3_1_13/a_109_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C16033 sky130_fd_sc_hd__or3b_2_0/a_176_21# sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# 0.00fF
C16034 sky130_fd_sc_hd__or3b_2_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# 0.00fF
C16035 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C16036 DOUT[9] DOUT[3] 0.03fF
C16037 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# VDD 0.06fF
C16038 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# sky130_fd_sc_hd__o221ai_1_0/a_109_47# 0.00fF
C16039 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# sky130_fd_sc_hd__o221ai_1_0/a_295_297# 0.00fF
C16040 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# sky130_fd_sc_hd__o221ai_1_0/a_213_123# 0.00fF
C16041 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# sky130_fd_sc_hd__o221ai_1_0/a_493_297# 0.00fF
C16042 sky130_fd_sc_hd__nor3_1_7/a_109_297# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C16043 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.00fF
C16044 sky130_fd_sc_hd__dfrtn_1_7/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C16045 sky130_fd_sc_hd__dfrtn_1_11/a_1462_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C16046 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C16047 sky130_fd_sc_hd__dfrtn_1_16/a_193_47# sky130_fd_sc_hd__inv_1_26/A 0.02fF
C16048 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C16049 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# VDD 0.00fF
C16050 sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C16051 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# DOUT[21] 0.00fF
C16052 DOUT[9] sky130_fd_sc_hd__inv_1_2/A 0.00fF
C16053 sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# sky130_fd_sc_hd__dfrtn_1_23/a_543_47# 0.00fF
C16054 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_6/a_193_47# 0.00fF
C16055 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C16056 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C16057 sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__inv_1_43/A 0.01fF
C16058 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__nor3_2_1/A 0.00fF
C16059 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# RESET_COUNTERn 0.00fF
C16060 sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C16061 sky130_fd_sc_hd__dfrtn_1_32/a_27_47# sky130_fd_sc_hd__inv_1_36/A 0.01fF
C16062 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C16063 DOUT[9] DOUT[5] 0.21fF
C16064 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# DOUT[3] 0.00fF
C16065 sky130_fd_sc_hd__nor3_2_3/B RESET_COUNTERn 2.82fF
C16066 sky130_fd_sc_hd__nor3_1_10/a_193_297# RESET_COUNTERn 0.00fF
C16067 sky130_fd_sc_hd__dfrtn_1_33/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C16068 sky130_fd_sc_hd__dfrtn_1_33/a_1270_413# VDD 0.00fF
C16069 sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# RESET_COUNTERn 0.02fF
C16070 sky130_fd_sc_hd__nor3_1_19/Y sky130_fd_sc_hd__o2111a_2_0/X 0.04fF
C16071 DOUT[1] sky130_fd_sc_hd__inv_1_39/A 0.83fF
C16072 sky130_fd_sc_hd__dfrtn_1_41/a_448_47# sky130_fd_sc_hd__inv_1_27/Y 0.00fF
C16073 sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C16074 sky130_fd_sc_hd__dfrtn_1_31/a_651_413# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C16075 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# DOUT[3] 0.00fF
C16076 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__or3_1_0/X 0.01fF
C16077 sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__dfrtn_1_9/a_27_47# -0.01fF
C16078 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__nor3_1_2/a_193_297# 0.00fF
C16079 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__nor3_1_19/Y 0.01fF
C16080 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# VDD 0.10fF
C16081 sky130_fd_sc_hd__dfrtn_1_20/a_1270_413# sky130_fd_sc_hd__inv_1_35/A 0.00fF
C16082 DOUT[4] sky130_fd_sc_hd__dfrtn_1_31/a_639_47# 0.00fF
C16083 sky130_fd_sc_hd__dfrtn_1_29/a_805_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C16084 sky130_fd_sc_hd__dfrtn_1_30/a_448_47# sky130_fd_sc_hd__dfrtn_1_31/a_448_47# 0.00fF
C16085 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# DOUT[14] 0.00fF
C16086 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C16087 sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# sky130_fd_sc_hd__inv_1_11/A 0.03fF
C16088 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C16089 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# sky130_fd_sc_hd__inv_1_15/A 0.03fF
C16090 sky130_fd_sc_hd__or2_2_0/X sky130_fd_sc_hd__dfrtn_1_17/a_805_47# 0.00fF
C16091 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# HEADER_0/a_508_138# 0.00fF
C16092 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__or2_2_0/B 0.02fF
C16093 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__nor3_2_3/C 0.05fF
C16094 sky130_fd_sc_hd__o211a_1_1/a_215_47# sky130_fd_sc_hd__dfrtn_1_17/a_639_47# 0.00fF
C16095 DOUT[13] sky130_fd_sc_hd__dfrtn_1_36/a_761_289# 0.00fF
C16096 sky130_fd_sc_hd__dfrtn_1_0/a_543_47# DOUT[17] 0.01fF
C16097 sky130_fd_sc_hd__dfrtn_1_34/a_805_47# SEL_CONV_TIME[1] 0.00fF
C16098 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# DOUT[6] 0.00fF
C16099 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# DOUT[20] 0.00fF
C16100 sky130_fd_sc_hd__dfrtn_1_24/a_1270_413# sky130_fd_sc_hd__dfrtn_1_29/a_27_47# 0.00fF
C16101 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# sky130_fd_sc_hd__dfrtn_1_29/a_448_47# 0.00fF
C16102 sky130_fd_sc_hd__dfrtn_1_24/a_651_413# sky130_fd_sc_hd__dfrtn_1_29/a_193_47# 0.00fF
C16103 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# 0.00fF
C16104 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_29/a_651_413# 0.00fF
C16105 sky130_fd_sc_hd__dfrtn_1_24/a_448_47# sky130_fd_sc_hd__dfrtn_1_29/a_761_289# 0.00fF
C16106 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__inv_1_28/A 0.01fF
C16107 sky130_fd_sc_hd__inv_1_38/A DOUT[21] 0.00fF
C16108 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C16109 sky130_fd_sc_hd__nand3b_1_1/a_53_93# RESET_COUNTERn 0.01fF
C16110 sky130_fd_sc_hd__nor3_1_5/a_193_297# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C16111 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# RESET_COUNTERn 0.06fF
C16112 sky130_fd_sc_hd__or3_1_0/a_29_53# RESET_COUNTERn 0.00fF
C16113 sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C16114 sky130_fd_sc_hd__dfrtn_1_38/a_448_47# VDD 0.04fF
C16115 sky130_fd_sc_hd__inv_1_31/A SEL_CONV_TIME[0] 0.24fF
C16116 sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# sky130_fd_sc_hd__inv_1_45/A 0.00fF
C16117 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C16118 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# 0.00fF
C16119 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_11/a_1217_47# 0.00fF
C16120 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_1462_47# 0.00fF
C16121 sky130_fd_sc_hd__dfrtn_1_10/a_805_47# sky130_fd_sc_hd__dfrtn_1_11/a_761_289# 0.00fF
C16122 sky130_fd_sc_hd__dfrtn_1_10/a_1270_413# sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# 0.00fF
C16123 sky130_fd_sc_hd__nor3_2_3/a_27_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C16124 sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# DOUT[15] 0.00fF
C16125 sky130_fd_sc_hd__nor3_1_4/a_109_297# DOUT[19] 0.00fF
C16126 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# 0.00fF
C16127 sky130_fd_sc_hd__inv_1_45/A DOUT[2] 0.00fF
C16128 sky130_fd_sc_hd__nor3_1_9/a_193_297# RESET_COUNTERn 0.00fF
C16129 sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C16130 sky130_fd_sc_hd__inv_1_33/Y DOUT[2] 0.25fF
C16131 sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# 0.00fF
C16132 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_17/a_1462_47# 0.00fF
C16133 sky130_fd_sc_hd__dfrtp_1_2/a_805_47# sky130_fd_sc_hd__dfrtn_1_17/a_651_413# 0.00fF
C16134 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# sky130_fd_sc_hd__dfrtn_1_17/a_805_47# 0.00fF
C16135 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__dfrtn_1_34/a_761_289# 0.00fF
C16136 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C16137 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__dfrtn_1_37/a_651_413# -0.00fF
C16138 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# 0.00fF
C16139 sky130_fd_sc_hd__dfrtn_1_28/a_639_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C16140 sky130_fd_sc_hd__dfrtn_1_26/a_448_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C16141 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C16142 sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# VDD 0.00fF
C16143 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# DOUT[14] 0.00fF
C16144 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# sky130_fd_sc_hd__dfrtn_1_41/a_761_289# -0.00fF
C16145 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C16146 sky130_fd_sc_hd__dfrtn_1_34/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C16147 sky130_fd_sc_hd__dfrtn_1_34/a_639_47# VDD 0.00fF
C16148 sky130_fd_sc_hd__dfrtn_1_3/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C16149 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__dfrtn_1_8/a_543_47# 0.00fF
C16150 sky130_fd_sc_hd__dfrtn_1_23/a_1270_413# sky130_fd_sc_hd__inv_1_40/Y 0.00fF
C16151 SLC_0/a_438_293# DOUT[15] 0.00fF
C16152 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# sky130_fd_sc_hd__inv_1_2/Y 0.01fF
C16153 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_3/a_448_47# -0.00fF
C16154 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# -0.00fF
C16155 sky130_fd_sc_hd__o221ai_1_0/a_109_47# SEL_CONV_TIME[0] 0.00fF
C16156 sky130_fd_sc_hd__nor3_1_13/a_193_297# sky130_fd_sc_hd__inv_1_9/Y 0.00fF
C16157 sky130_fd_sc_hd__dfrtn_1_25/a_1217_47# DOUT[21] 0.00fF
C16158 sky130_fd_sc_hd__dfrtn_1_25/a_448_47# RESET_COUNTERn 0.00fF
C16159 sky130_fd_sc_hd__dfrtp_1_3/a_761_289# sky130_fd_sc_hd__or2_2_0/X 0.01fF
C16160 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C16161 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# sky130_fd_sc_hd__or2_2_0/a_121_297# 0.00fF
C16162 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_5/Y 0.04fF
C16163 sky130_fd_sc_hd__inv_1_33/A SEL_CONV_TIME[0] 0.13fF
C16164 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# sky130_fd_sc_hd__inv_1_32/Y 0.00fF
C16165 sky130_fd_sc_hd__dfrtn_1_32/a_1217_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C16166 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# sky130_fd_sc_hd__inv_1_13/Y 0.00fF
C16167 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C16168 sky130_fd_sc_hd__inv_1_11/Y DOUT[21] -0.01fF
C16169 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# sky130_fd_sc_hd__or3b_2_0/X 0.00fF
C16170 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# sky130_fd_sc_hd__o211a_1_1/a_215_47# 0.00fF
C16171 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__o211a_1_1/a_510_47# 0.00fF
C16172 sky130_fd_sc_hd__dfrtp_1_3/a_543_47# sky130_fd_sc_hd__o211a_1_1/a_79_21# 0.00fF
C16173 DOUT[9] DOUT[20] 0.01fF
C16174 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# DOUT[15] 0.00fF
C16175 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# 0.03fF
C16176 DOUT[4] sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# 0.00fF
C16177 sky130_fd_sc_hd__nor3_1_8/a_109_297# DOUT[3] 0.00fF
C16178 sky130_fd_sc_hd__inv_1_47/A sky130_fd_sc_hd__inv_1_44/Y 0.01fF
C16179 sky130_fd_sc_hd__inv_1_17/A outb 0.00fF
C16180 sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C16181 sky130_fd_sc_hd__dfrtn_1_7/a_639_47# HEADER_0/a_508_138# 0.00fF
C16182 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_761_289# 0.00fF
C16183 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C16184 sky130_fd_sc_hd__dfrtn_1_28/a_543_47# SEL_CONV_TIME[1] 0.00fF
C16185 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C16186 sky130_fd_sc_hd__dfrtn_1_40/a_1462_47# VDD 0.00fF
C16187 sky130_fd_sc_hd__mux4_2_0/a_872_316# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C16188 sky130_fd_sc_hd__dfrtn_1_42/a_651_413# RESET_COUNTERn 0.00fF
C16189 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# SEL_CONV_TIME[3] 0.00fF
C16190 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__o311a_1_0/a_81_21# 0.00fF
C16191 sky130_fd_sc_hd__mux4_2_0/a_27_47# sky130_fd_sc_hd__o311a_1_0/a_585_47# 0.00fF
C16192 sky130_fd_sc_hd__nor3_2_3/B SEL_CONV_TIME[3] 0.03fF
C16193 sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C16194 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C16195 sky130_fd_sc_hd__inv_1_7/Y sky130_fd_sc_hd__nor3_2_3/B 0.58fF
C16196 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_10/a_651_413# 0.00fF
C16197 sky130_fd_sc_hd__dfrtn_1_0/a_1217_47# sky130_fd_sc_hd__inv_1_15/A 0.00fF
C16198 sky130_fd_sc_hd__nor3_1_10/a_193_297# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C16199 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__or3_1_0/C 0.02fF
C16200 sky130_fd_sc_hd__mux4_2_0/a_288_47# sky130_fd_sc_hd__mux4_2_0/a_372_413# -0.00fF
C16201 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtp_1_3/a_1108_47# 0.00fF
C16202 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# sky130_fd_sc_hd__dfrtp_1_3/a_639_47# 0.00fF
C16203 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# sky130_fd_sc_hd__dfrtp_1_3/a_448_47# 0.00fF
C16204 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C16205 sky130_fd_sc_hd__dfrtp_1_2/a_639_47# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.00fF
C16206 sky130_fd_sc_hd__nor2_1_0/a_109_297# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C16207 sky130_fd_sc_hd__o2111a_2_0/a_458_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C16208 sky130_fd_sc_hd__nor3_1_2/a_109_297# DOUT[18] 0.00fF
C16209 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# RESET_COUNTERn 0.00fF
C16210 sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# sky130_fd_sc_hd__inv_1_28/A 0.00fF
C16211 sky130_fd_sc_hd__inv_1_37/A sky130_fd_sc_hd__inv_1_13/A 0.12fF
C16212 sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# RESET_COUNTERn 0.00fF
C16213 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# SEL_CONV_TIME[0] 0.00fF
C16214 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C16215 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__nor3_1_3/a_193_297# 0.00fF
C16216 SLC_0/a_1235_416# RESET_COUNTERn 0.00fF
C16217 sky130_fd_sc_hd__nor3_1_10/a_109_297# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C16218 sky130_fd_sc_hd__dfrtn_1_31/a_448_47# sky130_fd_sc_hd__inv_1_49/A 0.00fF
C16219 DOUT[13] sky130_fd_sc_hd__dfrtn_1_31/a_1283_21# 0.00fF
C16220 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_761_289# 0.00fF
C16221 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_193_47# 0.00fF
C16222 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# SEL_CONV_TIME[2] 0.02fF
C16223 SLC_0/a_264_22# lc_out 0.02fF
C16224 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# 0.00fF
C16225 sky130_fd_sc_hd__dfrtn_1_28/a_761_289# VDD 0.06fF
C16226 sky130_fd_sc_hd__nand3b_1_1/a_53_93# SEL_CONV_TIME[3] 0.00fF
C16227 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_11/a_543_47# -0.00fF
C16228 sky130_fd_sc_hd__or3_1_0/a_29_53# SEL_CONV_TIME[3] 0.00fF
C16229 SEL_CONV_TIME[2] sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C16230 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# sky130_fd_sc_hd__o2111a_2_0/X 0.00fF
C16231 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__inv_1_7/Y 0.08fF
C16232 sky130_fd_sc_hd__dfrtn_1_14/a_651_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C16233 sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# sky130_fd_sc_hd__nor3_2_3/B 0.03fF
C16234 sky130_fd_sc_hd__dfrtn_1_14/a_639_47# VDD 0.00fF
C16235 sky130_fd_sc_hd__dfrtn_1_12/a_761_289# sky130_fd_sc_hd__dfrtn_1_0/a_1462_47# 0.00fF
C16236 sky130_fd_sc_hd__dfrtn_1_12/a_1462_47# sky130_fd_sc_hd__dfrtn_1_0/a_761_289# 0.00fF
C16237 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# sky130_fd_sc_hd__dfrtn_1_0/a_805_47# 0.00fF
C16238 sky130_fd_sc_hd__dfrtn_1_12/a_805_47# sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# 0.00fF
C16239 sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# sky130_fd_sc_hd__inv_1_2/Y 0.01fF
C16240 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_0/a_1270_413# 0.00fF
C16241 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__dfrtn_1_29/a_543_47# 0.00fF
C16242 sky130_fd_sc_hd__dfrtp_1_0/a_639_47# RESET_COUNTERn 0.00fF
C16243 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C16244 sky130_fd_sc_hd__dfrtn_1_41/a_1270_413# sky130_fd_sc_hd__inv_1_45/Y 0.00fF
C16245 DOUT[0] RESET_COUNTERn 0.00fF
C16246 sky130_fd_sc_hd__mux4_1_0/a_247_21# SEL_CONV_TIME[1] 0.00fF
C16247 sky130_fd_sc_hd__or3_1_0/X sky130_fd_sc_hd__inv_1_48/Y 0.08fF
C16248 sky130_fd_sc_hd__o221ai_1_0/a_493_297# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C16249 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__inv_1_41/Y 0.00fF
C16250 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# lc_out 0.00fF
C16251 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C16252 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C16253 lc_out DOUT[10] 0.03fF
C16254 sky130_fd_sc_hd__inv_1_2/Y DOUT[7] 0.00fF
C16255 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C16256 sky130_fd_sc_hd__nor3_1_14/a_193_297# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C16257 sky130_fd_sc_hd__dfrtn_1_24/a_651_413# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C16258 sky130_fd_sc_hd__dfrtn_1_39/a_805_47# RESET_COUNTERn 0.00fF
C16259 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# VDD 0.18fF
C16260 sky130_fd_sc_hd__dfrtn_1_22/a_1270_413# sky130_fd_sc_hd__inv_1_39/Y 0.00fF
C16261 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__inv_1_13/A 0.02fF
C16262 sky130_fd_sc_hd__dfrtn_1_42/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C16263 sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# DOUT[21] 0.01fF
C16264 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# sky130_fd_sc_hd__inv_1_42/A 0.01fF
C16265 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__nor3_1_3/a_193_297# 0.00fF
C16266 sky130_fd_sc_hd__nor3_1_16/a_193_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C16267 sky130_fd_sc_hd__dfrtn_1_18/a_805_47# RESET_COUNTERn 0.00fF
C16268 sky130_fd_sc_hd__or2b_1_0/a_27_53# sky130_fd_sc_hd__o2111a_2_0/a_80_21# 0.00fF
C16269 sky130_fd_sc_hd__or2b_1_0/a_219_297# sky130_fd_sc_hd__o2111a_2_0/a_674_297# 0.00fF
C16270 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C16271 sky130_fd_sc_hd__nor3_2_3/C sky130_fd_sc_hd__mux4_1_0/X 0.20fF
C16272 sky130_fd_sc_hd__or3_1_0/a_183_297# sky130_fd_sc_hd__dfrtn_1_25/a_761_289# 0.00fF
C16273 sky130_fd_sc_hd__or3_1_0/a_111_297# sky130_fd_sc_hd__dfrtn_1_25/a_543_47# 0.00fF
C16274 sky130_fd_sc_hd__dfrtn_1_20/a_543_47# sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# 0.00fF
C16275 DOUT[1] sky130_fd_sc_hd__dfrtn_1_36/a_27_47# 0.00fF
C16276 HEADER_0/a_508_138# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C16277 sky130_fd_sc_hd__dfrtn_1_23/a_761_289# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C16278 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C16279 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_26/a_193_47# 0.00fF
C16280 sky130_fd_sc_hd__dfrtn_1_22/a_761_289# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C16281 sky130_fd_sc_hd__dfrtn_1_4/a_639_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C16282 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# sky130_fd_sc_hd__dfrtn_1_42/a_193_47# -0.28fF
C16283 sky130_fd_sc_hd__dfrtn_1_25/a_448_47# SEL_CONV_TIME[3] 0.00fF
C16284 sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# SEL_CONV_TIME[0] 0.04fF
C16285 sky130_fd_sc_hd__dfrtn_1_3/a_639_47# sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# 0.00fF
C16286 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# 0.00fF
C16287 sky130_fd_sc_hd__mux4_1_0/a_193_413# VDD 0.01fF
C16288 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C16289 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# DOUT[3] 0.00fF
C16290 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C16291 SLC_0/a_264_22# sky130_fd_sc_hd__nor3_2_3/B 0.17fF
C16292 sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# VDD 0.07fF
C16293 sky130_fd_sc_hd__mux4_2_0/a_1281_47# sky130_fd_sc_hd__o311a_1_0/a_266_47# 0.00fF
C16294 sky130_fd_sc_hd__dfrtn_1_9/a_651_413# RESET_COUNTERn 0.01fF
C16295 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# sky130_fd_sc_hd__dfrtn_1_15/a_27_47# 0.00fF
C16296 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_761_289# 0.00fF
C16297 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_543_47# 0.00fF
C16298 sky130_fd_sc_hd__mux4_2_0/a_788_316# sky130_fd_sc_hd__mux4_2_0/a_1281_47# -0.00fF
C16299 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# DOUT[23] 0.00fF
C16300 sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C16301 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C16302 sky130_fd_sc_hd__dfrtn_1_19/a_448_47# RESET_COUNTERn 0.01fF
C16303 CLK_REF sky130_fd_sc_hd__dfrtn_1_17/a_805_47# 0.00fF
C16304 sky130_fd_sc_hd__nor3_1_8/a_109_297# DOUT[20] 0.00fF
C16305 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__inv_1_2/A 0.00fF
C16306 sky130_fd_sc_hd__o311a_1_0/a_266_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C16307 sky130_fd_sc_hd__dfrtn_1_41/a_805_47# sky130_fd_sc_hd__inv_1_43/A 0.00fF
C16308 sky130_fd_sc_hd__mux4_2_0/a_872_316# sky130_fd_sc_hd__inv_1_32/A 0.00fF
C16309 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__inv_1_49/A 0.01fF
C16310 sky130_fd_sc_hd__nand2_1_1/Y SEL_CONV_TIME[3] 0.02fF
C16311 sky130_fd_sc_hd__mux4_2_0/a_288_47# sky130_fd_sc_hd__inv_1_44/Y 0.00fF
C16312 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_761_289# -0.00fF
C16313 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_543_47# -0.00fF
C16314 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C16315 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# sky130_fd_sc_hd__dfrtn_1_4/a_543_47# 0.00fF
C16316 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_4/a_761_289# 0.00fF
C16317 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_4/a_448_47# 0.00fF
C16318 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_4/a_193_47# 0.00fF
C16319 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# sky130_fd_sc_hd__dfrtn_1_4/a_27_47# 0.00fF
C16320 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C16321 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C16322 sky130_fd_sc_hd__nor3_2_3/B DOUT[10] 0.03fF
C16323 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# sky130_fd_sc_hd__conb_1_0/LO 0.00fF
C16324 sky130_fd_sc_hd__dfrtn_1_37/a_639_47# sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# 0.00fF
C16325 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_1462_47# 0.00fF
C16326 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# 0.00fF
C16327 sky130_fd_sc_hd__nor3_1_2/a_193_297# RESET_COUNTERn 0.00fF
C16328 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C16329 sky130_fd_sc_hd__dfrtn_1_27/a_543_47# sky130_fd_sc_hd__inv_1_43/A 0.01fF
C16330 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__inv_1_5/A 0.00fF
C16331 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C16332 SEL_CONV_TIME[0] sky130_fd_sc_hd__o2111a_2_0/X 0.13fF
C16333 SEL_CONV_TIME[1] sky130_fd_sc_hd__inv_1_44/A 0.32fF
C16334 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_37/a_1270_413# 0.00fF
C16335 sky130_fd_sc_hd__dfrtn_1_21/a_1270_413# DOUT[2] 0.00fF
C16336 DOUT[23] sky130_fd_sc_hd__inv_1_40/Y 0.00fF
C16337 sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C16338 sky130_fd_sc_hd__dfrtn_1_9/a_639_47# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C16339 sky130_fd_sc_hd__dfrtn_1_0/a_448_47# VDD 0.01fF
C16340 sky130_fd_sc_hd__dfrtn_1_35/a_761_289# VDD 0.05fF
C16341 sky130_fd_sc_hd__dfrtn_1_12/a_761_289# sky130_fd_sc_hd__inv_1_15/A 0.03fF
C16342 sky130_fd_sc_hd__nor3_1_13/a_193_297# sky130_fd_sc_hd__dfrtn_1_8/a_193_47# 0.00fF
C16343 sky130_fd_sc_hd__dfrtn_1_11/a_639_47# sky130_fd_sc_hd__inv_1_37/A 0.00fF
C16344 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__inv_1_14/A 0.00fF
C16345 sky130_fd_sc_hd__mux4_2_0/X SEL_CONV_TIME[0] 0.12fF
C16346 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# DOUT[17] 0.00fF
C16347 sky130_fd_sc_hd__nor3_1_3/a_193_297# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C16348 sky130_fd_sc_hd__nor3_1_2/a_109_297# DOUT[22] 0.00fF
C16349 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_38/a_805_47# 0.00fF
C16350 sky130_fd_sc_hd__nand3b_1_1/Y sky130_fd_sc_hd__inv_1_41/Y 0.01fF
C16351 sky130_fd_sc_hd__nand2_1_1/Y SEL_CONV_TIME[2] 0.08fF
C16352 sky130_fd_sc_hd__dfrtn_1_27/a_193_47# sky130_fd_sc_hd__or3_1_0/C 0.48fF
C16353 sky130_fd_sc_hd__inv_1_29/Y sky130_fd_sc_hd__dfrtp_1_1/D 0.00fF
C16354 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# SEL_CONV_TIME[0] 0.02fF
C16355 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C16356 VDD sky130_fd_sc_hd__inv_1_8/Y 0.79fF
C16357 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# 0.00fF
C16358 sky130_fd_sc_hd__dfrtn_1_23/a_543_47# sky130_fd_sc_hd__inv_1_36/A 0.00fF
C16359 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# sky130_fd_sc_hd__inv_1_6/A 0.00fF
C16360 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_30/a_27_47# 0.00fF
C16361 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_24/a_761_289# 0.00fF
C16362 sky130_fd_sc_hd__dfrtn_1_20/a_1217_47# VDD 0.00fF
C16363 sky130_fd_sc_hd__dfrtn_1_24/a_805_47# RESET_COUNTERn 0.00fF
C16364 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_543_47# -0.00fF
C16365 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_761_289# -0.00fF
C16366 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# RESET_COUNTERn 0.03fF
C16367 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# sky130_fd_sc_hd__inv_1_26/A 0.01fF
C16368 sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C16369 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# SEL_CONV_TIME[1] 0.00fF
C16370 CLK_REF sky130_fd_sc_hd__dfrtp_1_3/a_761_289# 0.01fF
C16371 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# 0.01fF
C16372 DOUT[1] sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# 0.00fF
C16373 DOUT[4] sky130_fd_sc_hd__o311a_1_0/A3 0.02fF
C16374 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_4/a_1270_413# 0.00fF
C16375 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# -0.00fF
C16376 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# -0.00fF
C16377 sky130_fd_sc_hd__dfrtn_1_16/a_1270_413# DOUT[2] 0.00fF
C16378 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# sky130_fd_sc_hd__dfrtn_1_13/a_543_47# 0.00fF
C16379 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# 0.00fF
C16380 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# 0.00fF
C16381 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# sky130_fd_sc_hd__dfrtn_1_13/a_27_47# 0.00fF
C16382 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# sky130_fd_sc_hd__dfrtn_1_13/a_448_47# 0.00fF
C16383 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# VIN 0.07fF
C16384 DOUT[9] sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C16385 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# sky130_fd_sc_hd__inv_1_5/Y 0.01fF
C16386 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# DOUT[11] 0.00fF
C16387 sky130_fd_sc_hd__nor3_1_17/a_109_297# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C16388 sky130_fd_sc_hd__inv_1_47/Y DOUT[21] 0.20fF
C16389 sky130_fd_sc_hd__dfrtp_1_0/a_761_289# sky130_fd_sc_hd__dfrtp_1_0/a_543_47# -0.00fF
C16390 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# sky130_fd_sc_hd__dfrtp_1_0/a_1283_21# -0.00fF
C16391 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C16392 sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C16393 sky130_fd_sc_hd__mux4_1_0/a_834_97# VDD 0.01fF
C16394 sky130_fd_sc_hd__dfrtn_1_37/a_1270_413# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C16395 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# sky130_fd_sc_hd__inv_1_4/Y 0.01fF
C16396 sky130_fd_sc_hd__o211a_1_0/a_510_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C16397 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtn_1_19/a_639_47# 0.00fF
C16398 sky130_fd_sc_hd__dfrtn_1_11/a_639_47# sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# 0.00fF
C16399 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# 0.00fF
C16400 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# VIN 0.02fF
C16401 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# sky130_fd_sc_hd__inv_1_51/Y 0.00fF
C16402 sky130_fd_sc_hd__dfrtp_1_0/a_1462_47# DOUT[23] 0.00fF
C16403 sky130_fd_sc_hd__nor3_1_7/a_193_297# sky130_fd_sc_hd__inv_1_6/Y 0.00fF
C16404 sky130_fd_sc_hd__inv_1_33/Y sky130_fd_sc_hd__inv_1_30/Y 0.01fF
C16405 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# sky130_fd_sc_hd__dfrtn_1_27/a_805_47# -0.00fF
C16406 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# sky130_fd_sc_hd__inv_1_3/Y 0.01fF
C16407 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__inv_1_48/Y 0.01fF
C16408 sky130_fd_sc_hd__nor3_1_11/a_109_297# sky130_fd_sc_hd__inv_1_3/A 0.00fF
C16409 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C16410 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# RESET_COUNTERn 0.01fF
C16411 sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C16412 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_11/a_639_47# 0.00fF
C16413 sky130_fd_sc_hd__dfrtn_1_38/a_1270_413# SEL_CONV_TIME[0] 0.00fF
C16414 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# VDD 0.13fF
C16415 sky130_fd_sc_hd__nor3_2_0/a_281_297# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C16416 DOUT[4] sky130_fd_sc_hd__nor3_2_0/a_281_297# 0.01fF
C16417 sky130_fd_sc_hd__inv_1_37/A DOUT[12] 0.03fF
C16418 sky130_fd_sc_hd__inv_1_1/Y DOUT[11] 0.04fF
C16419 sky130_fd_sc_hd__or3_1_0/X sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C16420 sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C16421 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# DOUT[20] 0.00fF
C16422 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# RESET_COUNTERn 0.00fF
C16423 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__dfrtn_1_4/a_448_47# 0.00fF
C16424 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# 0.00fF
C16425 sky130_fd_sc_hd__dfrtn_1_39/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_448_47# -0.00fF
C16426 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_651_413# -0.00fF
C16427 sky130_fd_sc_hd__dfrtn_1_39/a_805_47# SEL_CONV_TIME[2] 0.00fF
C16428 sky130_fd_sc_hd__inv_1_47/Y sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C16429 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_39/a_761_289# 0.00fF
C16430 sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# sky130_fd_sc_hd__inv_1_35/A 0.01fF
C16431 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__inv_1_45/A 0.00fF
C16432 sky130_fd_sc_hd__dfrtn_1_39/a_543_47# sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# 0.00fF
C16433 DOUT[1] sky130_fd_sc_hd__dfrtn_1_32/a_651_413# 0.00fF
C16434 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__dfrtn_1_14/a_193_47# 0.00fF
C16435 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__dfrtn_1_14/a_761_289# 0.00fF
C16436 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_30/a_193_47# 0.00fF
C16437 sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# RESET_COUNTERn 0.00fF
C16438 sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# DOUT[19] 0.00fF
C16439 sky130_fd_sc_hd__a221oi_4_0/a_471_297# sky130_fd_sc_hd__mux4_2_0/a_872_316# 0.00fF
C16440 sky130_fd_sc_hd__a221oi_4_0/a_27_297# sky130_fd_sc_hd__mux4_2_0/a_1060_369# 0.00fF
C16441 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C16442 sky130_fd_sc_hd__dfrtn_1_30/a_639_47# RESET_COUNTERn 0.00fF
C16443 sky130_fd_sc_hd__inv_1_31/A sky130_fd_sc_hd__dfrtn_1_18/a_761_289# 0.01fF
C16444 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__inv_1_8/Y 0.08fF
C16445 outb DOUT[21] 0.08fF
C16446 sky130_fd_sc_hd__nor3_1_11/a_109_297# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C16447 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C16448 sky130_fd_sc_hd__dfrtn_1_3/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# 0.00fF
C16449 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.00fF
C16450 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C16451 sky130_fd_sc_hd__dfrtn_1_18/a_27_47# sky130_fd_sc_hd__dfrtn_1_18/a_651_413# -0.00fF
C16452 sky130_fd_sc_hd__dfrtn_1_18/a_193_47# sky130_fd_sc_hd__dfrtn_1_18/a_448_47# -0.00fF
C16453 sky130_fd_sc_hd__mux4_2_0/a_1279_413# SEL_CONV_TIME[1] 0.00fF
C16454 DOUT[2] RESET_COUNTERn 0.14fF
C16455 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# DOUT[19] 0.00fF
C16456 sky130_fd_sc_hd__dfrtn_1_27/a_1462_47# sky130_fd_sc_hd__or3_1_0/C 0.00fF
C16457 DOUT[19] DOUT[6] 0.03fF
C16458 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__or3_1_0/X 0.00fF
C16459 sky130_fd_sc_hd__dfrtn_1_34/a_1217_47# SEL_CONV_TIME[0] 0.00fF
C16460 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__or3_1_0/X 0.01fF
C16461 sky130_fd_sc_hd__dfrtn_1_17/a_193_47# sky130_fd_sc_hd__inv_1_34/Y 0.01fF
C16462 sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C16463 sky130_fd_sc_hd__inv_1_32/A SEL_CONV_TIME[1] 0.13fF
C16464 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C16465 sky130_fd_sc_hd__dfrtp_1_1/a_805_47# VDD 0.00fF
C16466 sky130_fd_sc_hd__inv_1_13/A DOUT[14] 0.01fF
C16467 sky130_fd_sc_hd__inv_1_50/A sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# 0.00fF
C16468 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__inv_1_12/A 0.00fF
C16469 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# sky130_fd_sc_hd__inv_1_47/A 0.01fF
C16470 sky130_fd_sc_hd__nor3_1_6/a_193_297# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C16471 sky130_fd_sc_hd__dfrtn_1_30/a_651_413# DONE 0.00fF
C16472 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C16473 sky130_fd_sc_hd__dfrtn_1_16/a_1108_47# sky130_fd_sc_hd__inv_1_25/A 0.00fF
C16474 sky130_fd_sc_hd__dfrtp_1_0/a_1270_413# SLC_0/a_919_243# 0.00fF
C16475 sky130_fd_sc_hd__dfrtp_1_0/a_639_47# SLC_0/a_264_22# 0.00fF
C16476 sky130_fd_sc_hd__dfrtp_1_0/a_805_47# SLC_0/a_438_293# 0.00fF
C16477 sky130_fd_sc_hd__inv_1_51/Y sky130_fd_sc_hd__inv_1_49/A 0.04fF
C16478 SLC_0/a_919_243# out 0.01fF
C16479 sky130_fd_sc_hd__dfrtp_1_0/a_1217_47# sky130_fd_sc_hd__inv_1_26/A 0.00fF
C16480 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C16481 sky130_fd_sc_hd__dfrtn_1_38/a_761_289# RESET_COUNTERn 0.05fF
C16482 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# DOUT[18] 0.01fF
C16483 VDD sky130_fd_sc_hd__inv_1_34/Y 0.18fF
C16484 DOUT[9] sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C16485 sky130_fd_sc_hd__nand3b_1_0/a_53_93# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C16486 sky130_fd_sc_hd__dfrtn_1_14/a_761_289# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C16487 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__nor3_1_5/a_109_297# 0.00fF
C16488 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C16489 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__dfrtn_1_24/a_1270_413# 0.00fF
C16490 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__o211a_1_1/X 0.02fF
C16491 sky130_fd_sc_hd__dfrtn_1_7/a_639_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C16492 sky130_fd_sc_hd__dfrtn_1_8/a_805_47# outb 0.00fF
C16493 sky130_fd_sc_hd__nor3_2_2/A sky130_fd_sc_hd__nor3_2_3/B 0.62fF
C16494 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# 0.03fF
C16495 sky130_fd_sc_hd__dfrtn_1_39/a_761_289# sky130_fd_sc_hd__inv_1_33/A 0.00fF
C16496 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_12/a_805_47# 0.00fF
C16497 sky130_fd_sc_hd__dfrtn_1_7/a_1217_47# VIN 0.00fF
C16498 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C16499 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C16500 sky130_fd_sc_hd__mux4_2_0/a_1060_369# VDD 0.00fF
C16501 sky130_fd_sc_hd__nor3_1_10/a_109_297# sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# 0.00fF
C16502 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__inv_1_7/Y 0.00fF
C16503 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# -0.27fF
C16504 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C16505 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# 0.00fF
C16506 sky130_fd_sc_hd__dfrtn_1_18/a_761_289# sky130_fd_sc_hd__inv_1_33/A 0.01fF
C16507 sky130_fd_sc_hd__dfrtn_1_27/a_448_47# SEL_CONV_TIME[1] 0.00fF
C16508 sky130_fd_sc_hd__inv_1_29/A sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# 0.02fF
C16509 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# RESET_COUNTERn 0.03fF
C16510 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# sky130_fd_sc_hd__inv_1_53/A 0.01fF
C16511 sky130_fd_sc_hd__dfrtp_1_1/a_639_47# sky130_fd_sc_hd__nor3_2_1/a_27_297# 0.00fF
C16512 sky130_fd_sc_hd__dfrtn_1_33/a_1108_47# sky130_fd_sc_hd__inv_1_43/Y 0.00fF
C16513 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C16514 sky130_fd_sc_hd__inv_1_53/A sky130_fd_sc_hd__nor3_2_3/B 0.21fF
C16515 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# sky130_fd_sc_hd__dfrtp_1_3/a_27_47# 0.01fF
C16516 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# sky130_fd_sc_hd__dfrtp_1_3/a_543_47# 0.00fF
C16517 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# sky130_fd_sc_hd__dfrtp_1_3/a_761_289# 0.01fF
C16518 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# sky130_fd_sc_hd__dfrtp_1_3/a_193_47# 0.00fF
C16519 sky130_fd_sc_hd__dfrtn_1_34/a_805_47# DOUT[21] 0.00fF
C16520 sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# RESET_COUNTERn 0.00fF
C16521 sky130_fd_sc_hd__dfrtn_1_33/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C16522 sky130_fd_sc_hd__dfrtn_1_35/a_1270_413# sky130_fd_sc_hd__inv_1_38/Y 0.00fF
C16523 sky130_fd_sc_hd__dfrtn_1_16/a_543_47# sky130_fd_sc_hd__nor3_2_3/A 0.01fF
C16524 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# VDD 0.01fF
C16525 sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C16526 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__or2b_1_0/X 0.00fF
C16527 sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# RESET_COUNTERn 0.00fF
C16528 sky130_fd_sc_hd__dfrtn_1_35/a_651_413# sky130_fd_sc_hd__inv_1_52/Y 0.00fF
C16529 sky130_fd_sc_hd__dfrtn_1_30/a_651_413# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C16530 sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# VDD 0.00fF
C16531 sky130_fd_sc_hd__nor3_1_8/a_193_297# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C16532 sky130_fd_sc_hd__dfrtn_1_3/a_1270_413# sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C16533 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# DOUT[2] 0.00fF
C16534 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_37/a_27_47# 0.00fF
C16535 sky130_fd_sc_hd__nor3_2_0/a_281_297# outb 0.00fF
C16536 sky130_fd_sc_hd__inv_1_37/A sky130_fd_sc_hd__nor3_2_3/C 0.07fF
C16537 sky130_fd_sc_hd__o211a_1_1/a_79_21# sky130_fd_sc_hd__dfrtp_1_1/D 0.00fF
C16538 sky130_fd_sc_hd__dfrtn_1_8/a_1108_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C16539 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.01fF
C16540 sky130_fd_sc_hd__inv_1_10/A sky130_fd_sc_hd__dfrtn_1_35/a_761_289# 0.00fF
C16541 sky130_fd_sc_hd__dfrtn_1_34/a_543_47# DONE 0.00fF
C16542 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__or3_1_0/X 0.00fF
C16543 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# 0.00fF
C16544 sky130_fd_sc_hd__dfrtn_1_28/a_1283_21# SEL_CONV_TIME[0] 0.00fF
C16545 sky130_fd_sc_hd__nand3b_1_0/Y sky130_fd_sc_hd__nand3b_1_0/a_232_47# 0.00fF
C16546 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__inv_1_31/A 0.00fF
C16547 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C16548 sky130_fd_sc_hd__dfrtn_1_27/a_543_47# sky130_fd_sc_hd__nor3_2_3/C 0.00fF
C16549 sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# sky130_fd_sc_hd__inv_1_8/Y 0.00fF
C16550 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C16551 sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# VDD 0.06fF
C16552 DOUT[23] sky130_fd_sc_hd__o211a_1_1/X 0.00fF
C16553 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# 0.00fF
C16554 sky130_fd_sc_hd__dfrtn_1_34/a_805_47# sky130_fd_sc_hd__o311a_1_0/A3 0.00fF
C16555 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# 0.00fF
C16556 sky130_fd_sc_hd__nor3_1_18/a_109_297# VDD 0.00fF
C16557 sky130_fd_sc_hd__nor3_1_9/a_193_297# sky130_fd_sc_hd__dfrtn_1_1/a_543_47# 0.00fF
C16558 sky130_fd_sc_hd__nor3_1_9/a_109_297# sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# 0.00fF
C16559 sky130_fd_sc_hd__dfrtn_1_40/a_1270_413# RESET_COUNTERn 0.00fF
C16560 sky130_fd_sc_hd__dfrtp_1_2/a_448_47# sky130_fd_sc_hd__dfrtp_1_1/D 0.00fF
C16561 sky130_fd_sc_hd__dfrtn_1_17/a_1462_47# sky130_fd_sc_hd__inv_1_34/Y 0.00fF
C16562 sky130_fd_sc_hd__nor3_1_6/a_109_297# sky130_fd_sc_hd__inv_1_7/A 0.00fF
C16563 sky130_fd_sc_hd__dfrtn_1_36/a_193_47# sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# -0.00fF
C16564 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# -0.00fF
C16565 sky130_fd_sc_hd__dfrtn_1_36/a_761_289# sky130_fd_sc_hd__dfrtn_1_36/a_543_47# -0.00fF
C16566 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# sky130_fd_sc_hd__inv_1_13/A 0.00fF
C16567 sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# sky130_fd_sc_hd__inv_1_47/A 0.00fF
C16568 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__inv_1_53/Y 0.00fF
C16569 sky130_fd_sc_hd__o2111a_2_0/a_674_297# RESET_COUNTERn 0.00fF
C16570 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# sky130_fd_sc_hd__inv_1_6/A 0.02fF
C16571 sky130_fd_sc_hd__conb_1_0/LO DOUT[15] 0.00fF
C16572 sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# sky130_fd_sc_hd__inv_1_11/Y 0.00fF
C16573 sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# sky130_fd_sc_hd__inv_1_43/Y 0.02fF
C16574 sky130_fd_sc_hd__nor3_2_3/B sky130_fd_sc_hd__inv_1_4/Y 0.44fF
C16575 sky130_fd_sc_hd__nor3_1_10/a_193_297# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C16576 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# DOUT[18] 0.00fF
C16577 sky130_fd_sc_hd__inv_1_42/Y sky130_fd_sc_hd__nor3_2_3/B 0.08fF
C16578 sky130_fd_sc_hd__dfrtn_1_26/a_761_289# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C16579 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# sky130_fd_sc_hd__nor3_2_3/C 0.01fF
C16580 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# VDD 0.00fF
C16581 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_5/a_651_413# 0.00fF
C16582 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# sky130_fd_sc_hd__dfrtn_1_5/a_639_47# 0.00fF
C16583 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# sky130_fd_sc_hd__dfrtn_1_5/a_27_47# 0.00fF
C16584 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__dfrtn_1_5/a_543_47# 0.00fF
C16585 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# sky130_fd_sc_hd__dfrtn_1_5/a_193_47# 0.00fF
C16586 sky130_fd_sc_hd__nor3_1_19/a_109_297# RESET_COUNTERn 0.00fF
C16587 sky130_fd_sc_hd__dfrtp_1_3/a_651_413# sky130_fd_sc_hd__or2_2_0/B 0.00fF
C16588 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__nor3_1_1/a_193_297# 0.00fF
C16589 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__o221ai_1_0/a_295_297# 0.00fF
C16590 sky130_fd_sc_hd__inv_1_45/A sky130_fd_sc_hd__dfrtn_1_27/a_193_47# 0.01fF
C16591 sky130_fd_sc_hd__a221oi_4_0/a_471_297# SEL_CONV_TIME[1] 0.01fF
C16592 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# sky130_fd_sc_hd__inv_1_44/A 0.00fF
C16593 sky130_fd_sc_hd__dfrtn_1_34/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.02fF
C16594 sky130_fd_sc_hd__dfrtn_1_12/a_1270_413# VDD 0.00fF
C16595 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_30/a_448_47# 0.00fF
C16596 sky130_fd_sc_hd__dfrtp_1_2/a_805_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C16597 sky130_fd_sc_hd__dfrtn_1_17/a_639_47# sky130_fd_sc_hd__inv_1_28/Y 0.00fF
C16598 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__nor3_2_3/C 0.50fF
C16599 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__dfrtn_1_1/a_761_289# 0.00fF
C16600 sky130_fd_sc_hd__inv_1_8/Y DOUT[3] 0.00fF
C16601 sky130_fd_sc_hd__dfrtn_1_28/a_543_47# DOUT[21] 0.01fF
C16602 sky130_fd_sc_hd__dfrtn_1_14/a_761_289# sky130_fd_sc_hd__nor3_1_1/a_109_297# 0.00fF
C16603 sky130_fd_sc_hd__dfrtn_1_33/a_651_413# DOUT[23] 0.00fF
C16604 sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C16605 sky130_fd_sc_hd__dfrtn_1_0/a_448_47# DOUT[5] 0.00fF
C16606 sky130_fd_sc_hd__dfrtn_1_11/a_639_47# DOUT[14] 0.00fF
C16607 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# RESET_COUNTERn 0.01fF
C16608 sky130_fd_sc_hd__mux4_1_0/a_277_47# SEL_CONV_TIME[0] 0.01fF
C16609 sky130_fd_sc_hd__dfrtn_1_28/a_651_413# sky130_fd_sc_hd__inv_1_48/Y 0.00fF
C16610 sky130_fd_sc_hd__inv_1_30/A sky130_fd_sc_hd__inv_1_33/A 0.00fF
C16611 sky130_fd_sc_hd__dfrtn_1_42/a_651_413# sky130_fd_sc_hd__nor3_2_2/A 0.00fF
C16612 sky130_fd_sc_hd__or3b_2_0/B sky130_fd_sc_hd__dfrtn_1_34/a_1270_413# 0.00fF
C16613 sky130_fd_sc_hd__or3b_2_0/a_176_21# SEL_CONV_TIME[1] 0.02fF
C16614 sky130_fd_sc_hd__nor3_1_8/a_109_297# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C16615 sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# sky130_fd_sc_hd__dfrtp_1_3/a_761_289# 0.00fF
C16616 sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# sky130_fd_sc_hd__dfrtp_1_3/a_543_47# 0.00fF
C16617 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# sky130_fd_sc_hd__dfrtp_1_3/a_639_47# 0.00fF
C16618 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C16619 sky130_fd_sc_hd__dfrtn_1_20/a_448_47# sky130_fd_sc_hd__dfrtn_1_21/a_761_289# 0.00fF
C16620 sky130_fd_sc_hd__dfrtn_1_20/a_651_413# sky130_fd_sc_hd__dfrtn_1_21/a_1270_413# 0.00fF
C16621 sky130_fd_sc_hd__or3_1_0/a_29_53# sky130_fd_sc_hd__inv_1_42/Y 0.01fF
C16622 sky130_fd_sc_hd__dfrtn_1_36/a_1270_413# sky130_fd_sc_hd__inv_1_40/A 0.00fF
C16623 sky130_fd_sc_hd__dfrtn_1_4/a_761_289# VIN 0.00fF
C16624 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# DOUT[22] 0.00fF
C16625 DOUT[9] sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C16626 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# sky130_fd_sc_hd__dfrtn_1_37/a_639_47# 0.00fF
C16627 sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# sky130_fd_sc_hd__dfrtn_1_37/a_27_47# 0.00fF
C16628 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# sky130_fd_sc_hd__dfrtn_1_37/a_193_47# 0.00fF
C16629 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_37/a_805_47# 0.00fF
C16630 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# sky130_fd_sc_hd__inv_1_48/A 0.00fF
C16631 sky130_fd_sc_hd__nand3b_1_1/a_53_93# sky130_fd_sc_hd__dfrtn_1_34/a_543_47# 0.00fF
C16632 sky130_fd_sc_hd__nand3b_1_1/a_316_47# sky130_fd_sc_hd__dfrtn_1_34/a_193_47# 0.00fF
C16633 sky130_fd_sc_hd__nor3_1_1/a_193_297# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C16634 sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__inv_1_53/A 0.00fF
C16635 sky130_fd_sc_hd__a221oi_4_0/a_27_297# VDD 0.11fF
C16636 VDD sky130_fd_sc_hd__inv_1_40/A 0.37fF
C16637 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# sky130_fd_sc_hd__dfrtn_1_2/a_543_47# 0.00fF
C16638 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__dfrtn_1_2/a_761_289# 0.00fF
C16639 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# sky130_fd_sc_hd__dfrtn_1_2/a_193_47# 0.00fF
C16640 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# 0.00fF
C16641 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# sky130_fd_sc_hd__dfrtn_1_2/a_27_47# 0.00fF
C16642 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# sky130_fd_sc_hd__dfrtn_1_2/a_448_47# 0.00fF
C16643 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# 0.00fF
C16644 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__dfrtn_1_2/a_805_47# 0.00fF
C16645 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# 0.00fF
C16646 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# sky130_fd_sc_hd__dfrtn_1_2/a_639_47# 0.00fF
C16647 sky130_fd_sc_hd__inv_1_46/Y sky130_fd_sc_hd__dfrtn_1_25/a_761_289# 0.00fF
C16648 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# sky130_fd_sc_hd__nor3_2_0/A 0.00fF
C16649 sky130_fd_sc_hd__dfrtn_1_22/a_543_47# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C16650 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# sky130_fd_sc_hd__dfrtn_1_24/a_651_413# -0.00fF
C16651 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# sky130_fd_sc_hd__dfrtn_1_24/a_448_47# -0.00fF
C16652 sky130_fd_sc_hd__dfrtp_1_3/a_805_47# sky130_fd_sc_hd__or2_2_0/a_39_297# 0.00fF
C16653 DOUT[9] sky130_fd_sc_hd__dfrtn_1_5/a_805_47# 0.00fF
C16654 sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# sky130_fd_sc_hd__nor3_2_3/B 0.00fF
C16655 sky130_fd_sc_hd__dfrtn_1_39/a_651_413# sky130_fd_sc_hd__inv_1_31/Y 0.00fF
C16656 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# sky130_fd_sc_hd__dfrtn_1_17/a_761_289# -0.00fF
C16657 DOUT[1] sky130_fd_sc_hd__dfrtn_1_22/a_639_47# 0.00fF
C16658 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__dfrtn_1_34/a_761_289# 0.01fF
C16659 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# SEL_CONV_TIME[1] 0.01fF
C16660 DOUT[4] sky130_fd_sc_hd__o221ai_1_0/a_295_297# 0.00fF
C16661 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__inv_1_45/Y 0.01fF
C16662 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# DOUT[21] 0.00fF
C16663 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# RESET_COUNTERn -0.02fF
C16664 sky130_fd_sc_hd__inv_1_27/A sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# 0.02fF
C16665 DOUT[11] RESET_COUNTERn 0.03fF
C16666 sky130_fd_sc_hd__inv_1_34/A sky130_fd_sc_hd__dfrtn_1_19/a_761_289# 0.01fF
C16667 sky130_fd_sc_hd__dfrtn_1_26/a_651_413# DOUT[23] 0.00fF
C16668 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# DOUT[19] 0.01fF
C16669 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# DOUT[14] 0.00fF
C16670 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# sky130_fd_sc_hd__dfrtn_1_15/a_651_413# 0.00fF
C16671 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# 0.00fF
C16672 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# sky130_fd_sc_hd__dfrtn_1_15/a_761_289# 0.00fF
C16673 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# 0.00fF
C16674 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# 0.00fF
C16675 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# sky130_fd_sc_hd__dfrtn_1_15/a_193_47# 0.00fF
C16676 DOUT[12] DOUT[14] 0.02fF
C16677 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C16678 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# 0.00fF
C16679 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# sky130_fd_sc_hd__dfrtn_1_9/a_639_47# 0.00fF
C16680 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# sky130_fd_sc_hd__dfrtn_1_9/a_805_47# 0.00fF
C16681 sky130_fd_sc_hd__dfrtn_1_5/a_805_47# sky130_fd_sc_hd__dfrtn_1_9/a_27_47# 0.00fF
C16682 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C16683 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# sky130_fd_sc_hd__dfrtn_1_9/a_193_47# 0.00fF
C16684 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C16685 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# 0.00fF
C16686 sky130_fd_sc_hd__dfrtn_1_17/a_193_47# VDD 0.08fF
C16687 sky130_fd_sc_hd__dfrtn_1_25/a_448_47# sky130_fd_sc_hd__inv_1_42/Y 0.00fF
C16688 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__inv_1_54/Y 0.00fF
C16689 sky130_fd_sc_hd__dfrtn_1_14/a_651_413# sky130_fd_sc_hd__nor3_1_0/a_109_297# 0.00fF
C16690 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# sky130_fd_sc_hd__inv_1_8/A 0.00fF
C16691 sky130_fd_sc_hd__dfrtn_1_14/a_543_47# sky130_fd_sc_hd__nor3_2_3/B 0.01fF
C16692 sky130_fd_sc_hd__dfrtn_1_36/a_1270_413# VDD 0.00fF
C16693 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# 0.00fF
C16694 sky130_fd_sc_hd__a221oi_4_0/a_453_47# sky130_fd_sc_hd__nor3_1_19/Y 0.00fF
C16695 sky130_fd_sc_hd__dfrtn_1_40/a_1270_413# SEL_CONV_TIME[3] 0.00fF
C16696 sky130_fd_sc_hd__nor3_2_3/a_281_297# sky130_fd_sc_hd__dfrtn_1_42/a_761_289# 0.00fF
C16697 sky130_fd_sc_hd__nor3_2_3/a_27_297# sky130_fd_sc_hd__dfrtn_1_42/a_543_47# 0.00fF
C16698 sky130_fd_sc_hd__nor3_1_5/A sky130_fd_sc_hd__dfrtn_1_13/a_543_47# 0.00fF
C16699 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# sky130_fd_sc_hd__inv_1_2/Y 0.00fF
C16700 sky130_fd_sc_hd__dfrtn_1_0/a_805_47# sky130_fd_sc_hd__nor3_1_0/A 0.00fF
C16701 sky130_fd_sc_hd__dfrtn_1_17/a_1270_413# sky130_fd_sc_hd__or2_2_0/A 0.00fF
C16702 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# sky130_fd_sc_hd__inv_1_5/A 0.02fF
C16703 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# sky130_fd_sc_hd__inv_1_5/Y 0.00fF
C16704 sky130_fd_sc_hd__o2111a_2_0/a_674_297# SEL_CONV_TIME[3] 0.00fF
C16705 sky130_fd_sc_hd__o311a_1_0/a_81_21# sky130_fd_sc_hd__nand3b_1_1/Y 0.00fF
C16706 sky130_fd_sc_hd__inv_1_25/A DOUT[23] 0.00fF
C16707 sky130_fd_sc_hd__dfrtn_1_28/a_639_47# RESET_COUNTERn 0.00fF
C16708 sky130_fd_sc_hd__dfrtn_1_30/a_805_47# sky130_fd_sc_hd__inv_1_50/Y 0.00fF
C16709 sky130_fd_sc_hd__dfrtn_1_39/a_805_47# sky130_fd_sc_hd__inv_1_53/A 0.00fF
C16710 sky130_fd_sc_hd__dfrtn_1_0/a_761_289# RESET_COUNTERn 0.01fF
C16711 sky130_fd_sc_hd__dfrtn_1_35/a_543_47# DOUT[21] 0.00fF
C16712 sky130_fd_sc_hd__inv_1_52/A sky130_fd_sc_hd__inv_1_36/A 0.06fF
C16713 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# sky130_fd_sc_hd__inv_1_1/A 0.00fF
C16714 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# sky130_fd_sc_hd__or2b_1_0/X 0.01fF
C16715 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# sky130_fd_sc_hd__inv_1_39/A 0.00fF
C16716 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# sky130_fd_sc_hd__inv_1_4/Y 0.00fF
C16717 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# 0.00fF
C16718 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# 0.00fF
C16719 sky130_fd_sc_hd__inv_1_49/Y sky130_fd_sc_hd__dfrtn_1_30/a_761_289# 0.00fF
C16720 sky130_fd_sc_hd__dfrtn_1_40/a_1270_413# SEL_CONV_TIME[2] 0.00fF
C16721 sky130_fd_sc_hd__nor3_1_3/a_109_297# sky130_fd_sc_hd__nor3_1_4/A 0.00fF
C16722 sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# sky130_fd_sc_hd__dfrtn_1_36/a_1270_413# 0.00fF
C16723 sky130_fd_sc_hd__dfrtn_1_32/a_1270_413# sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# 0.00fF
C16724 sky130_fd_sc_hd__nor3_1_5/a_109_297# RESET_COUNTERn 0.00fF
C16725 sky130_fd_sc_hd__nand2_1_2/Y sky130_fd_sc_hd__inv_1_49/A 0.00fF
C16726 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# sky130_fd_sc_hd__inv_1_3/Y 0.00fF
C16727 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# sky130_fd_sc_hd__dfrtn_1_9/a_651_413# 0.00fF
C16728 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# sky130_fd_sc_hd__dfrtn_1_9/a_543_47# 0.00fF
C16729 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# sky130_fd_sc_hd__dfrtn_1_19/a_27_47# 0.00fF
C16730 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# sky130_fd_sc_hd__dfrtn_1_19/a_193_47# 0.00fF
C16731 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# DOUT[22] 0.00fF
C16732 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# sky130_fd_sc_hd__inv_1_31/A 0.15fF
C16733 DOUT[14] VSS 5.59fF
C16734 DOUT[18] VSS 2.85fF
C16735 DOUT[3] VSS 2.37fF
C16736 RESET_COUNTERn VSS 24.57fF
C16737 DOUT[8] VSS 4.74fF
C16738 DOUT[7] VSS 3.17fF
C16739 DOUT[6] VSS 2.78fF
C16740 DOUT[20] VSS 1.55fF
C16741 DOUT[21] VSS 3.04fF
C16742 SEL_CONV_TIME[3] VSS 1.92fF
C16743 DOUT[0] VSS 4.53fF
C16744 out VSS 8.92fF
C16745 DOUT[10] VSS 11.67fF
C16746 VIN VSS 166.17fF
C16747 DOUT[17] VSS 4.57fF
C16748 sky130_fd_sc_hd__nor3_1_0/A VSS 0.50fF
C16749 DOUT[1] VSS 4.64fF
C16750 sky130_fd_sc_hd__or3b_2_0/B VSS 0.72fF
C16751 DOUT[4] VSS 5.93fF
C16752 sky130_fd_sc_hd__inv_1_1/Y VSS 0.69fF
C16753 sky130_fd_sc_hd__nor3_1_5/A VSS 1.10fF
C16754 sky130_fd_sc_hd__inv_1_50/A VSS 0.44fF
C16755 sky130_fd_sc_hd__nand2_1_2/Y VSS 0.08fF
C16756 sky130_fd_sc_hd__inv_1_49/A VSS 2.47fF
C16757 sky130_fd_sc_hd__inv_1_51/Y VSS 0.46fF
C16758 sky130_fd_sc_hd__inv_1_8/A VSS 0.67fF
C16759 sky130_fd_sc_hd__inv_1_8/Y VSS 0.45fF
C16760 sky130_fd_sc_hd__inv_1_2/Y VSS 0.39fF
C16761 sky130_fd_sc_hd__inv_1_5/A VSS 0.41fF
C16762 sky130_fd_sc_hd__inv_1_13/A VSS 0.31fF
C16763 sky130_fd_sc_hd__inv_1_5/Y VSS 1.28fF
C16764 sky130_fd_sc_hd__inv_1_6/A VSS 1.09fF
C16765 sky130_fd_sc_hd__inv_1_4/Y VSS 0.41fF
C16766 sky130_fd_sc_hd__inv_1_6/Y VSS 0.33fF
C16767 sky130_fd_sc_hd__inv_1_12/A VSS 0.62fF
C16768 sky130_fd_sc_hd__inv_1_13/Y VSS 0.61fF
C16769 sky130_fd_sc_hd__nor3_1_4/A VSS 0.29fF
C16770 sky130_fd_sc_hd__inv_1_40/A VSS 0.62fF
C16771 sky130_fd_sc_hd__inv_1_38/Y VSS 0.91fF
C16772 sky130_fd_sc_hd__inv_1_40/Y VSS 1.11fF
C16773 sky130_fd_sc_hd__inv_1_3/A VSS 0.54fF
C16774 sky130_fd_sc_hd__nor3_2_3/B VSS 11.12fF
C16775 sky130_fd_sc_hd__inv_1_3/Y VSS 2.15fF
C16776 DOUT[19] VSS 8.14fF
C16777 sky130_fd_sc_hd__inv_1_39/Y VSS 0.40fF
C16778 sky130_fd_sc_hd__inv_1_43/A VSS 0.55fF
C16779 sky130_fd_sc_hd__inv_1_48/Y VSS 0.13fF
C16780 sky130_fd_sc_hd__inv_1_48/A VSS 1.18fF
C16781 sky130_fd_sc_hd__or3_1_0/C VSS 0.38fF
C16782 sky130_fd_sc_hd__o2111a_2_0/X VSS 0.27fF
C16783 sky130_fd_sc_hd__inv_1_44/A VSS 0.31fF
C16784 sky130_fd_sc_hd__inv_1_44/Y VSS 0.31fF
C16785 sky130_fd_sc_hd__o311a_1_0/A3 VSS 2.86fF
C16786 SEL_CONV_TIME[2] VSS 2.89fF
C16787 sky130_fd_sc_hd__inv_1_41/Y VSS 0.43fF
C16788 sky130_fd_sc_hd__mux4_1_0/X VSS 0.40fF
C16789 SEL_CONV_TIME[1] VSS 6.05fF
C16790 SEL_CONV_TIME[0] VSS 4.01fF
C16791 sky130_fd_sc_hd__inv_1_43/Y VSS 0.41fF
C16792 sky130_fd_sc_hd__inv_1_53/A VSS 1.01fF
C16793 sky130_fd_sc_hd__inv_1_53/Y VSS 0.29fF
C16794 sky130_fd_sc_hd__inv_1_32/Y VSS 0.27fF
C16795 sky130_fd_sc_hd__inv_1_33/A VSS 0.41fF
C16796 DOUT[2] VSS 5.34fF
C16797 sky130_fd_sc_hd__nor3_2_3/A VSS 1.02fF
C16798 sky130_fd_sc_hd__inv_1_23/A VSS 0.92fF
C16799 DOUT[12] VSS 4.54fF
C16800 lc_out VSS 3.62fF
C16801 sky130_fd_sc_hd__or2_2_0/A VSS 0.61fF
C16802 sky130_fd_sc_hd__inv_1_35/Y VSS 0.11fF
C16803 sky130_fd_sc_hd__inv_1_30/Y VSS 0.44fF
C16804 sky130_fd_sc_hd__o211a_1_0/X VSS 0.19fF
C16805 sky130_fd_sc_hd__dfrtp_1_1/D VSS 0.50fF
C16806 sky130_fd_sc_hd__o211a_1_1/X VSS 0.21fF
C16807 sky130_fd_sc_hd__inv_1_28/Y VSS 0.19fF
C16808 DOUT[15] VSS 3.53fF
C16809 DOUT[23] VSS 13.12fF
C16810 sky130_fd_sc_hd__inv_1_15/A VSS 2.31fF
C16811 sky130_fd_sc_hd__nor3_2_3/C VSS 15.25fF
C16812 DOUT[5] VSS 9.80fF
C16813 DOUT[22] VSS 2.87fF
C16814 sky130_fd_sc_hd__inv_1_7/A VSS 0.31fF
C16815 sky130_fd_sc_hd__inv_1_1/A VSS 3.95fF
C16816 DOUT[11] VSS 3.05fF
C16817 sky130_fd_sc_hd__nor3_2_0/A VSS 0.81fF
C16818 sky130_fd_sc_hd__inv_1_0/Y VSS 0.28fF
C16819 sky130_fd_sc_hd__inv_1_11/A VSS 0.23fF
C16820 sky130_fd_sc_hd__inv_1_11/Y VSS 1.83fF
C16821 en VSS 6.51fF
C16822 sky130_fd_sc_hd__inv_1_22/A VSS 0.36fF
C16823 sky130_fd_sc_hd__inv_1_19/A VSS 0.40fF
C16824 sky130_fd_sc_hd__inv_1_22/Y VSS 0.40fF
C16825 outb VSS 8.08fF
C16826 sky130_fd_sc_hd__inv_1_24/A VSS 0.25fF
C16827 sky130_fd_sc_hd__inv_1_17/A VSS 0.25fF
C16828 sky130_fd_sc_hd__inv_1_9/A VSS 1.74fF
C16829 sky130_fd_sc_hd__inv_1_9/Y VSS 0.53fF
C16830 sky130_fd_sc_hd__inv_1_36/Y VSS 0.59fF
C16831 sky130_fd_sc_hd__inv_1_36/A VSS 1.18fF
C16832 sky130_fd_sc_hd__inv_1_39/A VSS 0.60fF
C16833 sky130_fd_sc_hd__inv_1_52/Y VSS 0.54fF
C16834 sky130_fd_sc_hd__nor3_2_2/A VSS 0.43fF
C16835 sky130_fd_sc_hd__inv_1_25/A VSS 0.37fF
C16836 sky130_fd_sc_hd__inv_1_37/A VSS 2.17fF
C16837 sky130_fd_sc_hd__or2_2_0/B VSS 0.52fF
C16838 sky130_fd_sc_hd__inv_1_38/A VSS 0.47fF
C16839 DOUT[16] VSS 2.74fF
C16840 sky130_fd_sc_hd__inv_1_26/A VSS 0.36fF
C16841 sky130_fd_sc_hd__inv_1_29/Y VSS 0.13fF
C16842 sky130_fd_sc_hd__inv_1_42/A VSS 0.70fF
C16843 sky130_fd_sc_hd__or3_1_0/X VSS 0.14fF
C16844 sky130_fd_sc_hd__inv_1_28/A VSS 0.34fF
C16845 sky130_fd_sc_hd__inv_1_27/Y VSS 0.32fF
C16846 sky130_fd_sc_hd__inv_1_34/Y VSS 0.45fF
C16847 sky130_fd_sc_hd__inv_1_50/Y VSS 0.30fF
C16848 sky130_fd_sc_hd__or2b_1_0/X VSS 0.28fF
C16849 sky130_fd_sc_hd__nor3_1_19/Y VSS 0.14fF
C16850 sky130_fd_sc_hd__inv_1_35/A VSS 0.32fF
C16851 sky130_fd_sc_hd__nand3b_1_1/Y VSS 0.13fF
C16852 sky130_fd_sc_hd__nand2_1_1/Y VSS 0.26fF
C16853 sky130_fd_sc_hd__or3b_2_0/X VSS 0.16fF
C16854 DONE VSS 2.42fF
C16855 sky130_fd_sc_hd__inv_1_47/A VSS 0.53fF
C16856 sky130_fd_sc_hd__inv_1_31/Y VSS 0.10fF
C16857 sky130_fd_sc_hd__inv_1_32/A VSS 0.36fF
C16858 sky130_fd_sc_hd__nor3_1_5/a_193_297# VSS 0.00fF
C16859 sky130_fd_sc_hd__nor3_1_5/a_109_297# VSS 0.00fF
C16860 sky130_fd_sc_hd__dfrtn_1_9/a_1462_47# VSS 0.00fF
C16861 sky130_fd_sc_hd__dfrtn_1_9/a_1217_47# VSS 0.00fF
C16862 sky130_fd_sc_hd__dfrtn_1_9/a_805_47# VSS 0.00fF
C16863 sky130_fd_sc_hd__dfrtn_1_9/a_639_47# VSS 0.00fF
C16864 sky130_fd_sc_hd__dfrtn_1_9/a_1270_413# VSS 0.00fF
C16865 sky130_fd_sc_hd__dfrtn_1_9/a_651_413# VSS 0.01fF
C16866 sky130_fd_sc_hd__dfrtn_1_9/a_448_47# VSS 0.02fF
C16867 sky130_fd_sc_hd__dfrtn_1_9/a_1108_47# VSS 0.16fF
C16868 sky130_fd_sc_hd__dfrtn_1_9/a_1283_21# VSS 0.30fF
C16869 sky130_fd_sc_hd__dfrtn_1_9/a_543_47# VSS 0.16fF
C16870 sky130_fd_sc_hd__dfrtn_1_9/a_761_289# VSS 0.13fF
C16871 sky130_fd_sc_hd__dfrtn_1_9/a_193_47# VSS 0.23fF
C16872 sky130_fd_sc_hd__dfrtn_1_9/a_27_47# VSS 0.46fF
C16873 HEADER_0/a_508_138# VSS 0.13fF
C16874 VDD VSS 988.15fF
C16875 sky130_fd_sc_hd__inv_1_2/A VSS 1.93fF
C16876 sky130_fd_sc_hd__inv_1_42/Y VSS 0.46fF
C16877 sky130_fd_sc_hd__inv_1_7/Y VSS 0.21fF
C16878 sky130_fd_sc_hd__nor3_1_4/a_193_297# VSS 0.00fF
C16879 sky130_fd_sc_hd__nor3_1_4/a_109_297# VSS 0.00fF
C16880 sky130_fd_sc_hd__dfrtn_1_8/a_1462_47# VSS 0.01fF
C16881 sky130_fd_sc_hd__dfrtn_1_8/a_1217_47# VSS 0.00fF
C16882 sky130_fd_sc_hd__dfrtn_1_8/a_805_47# VSS 0.00fF
C16883 sky130_fd_sc_hd__dfrtn_1_8/a_639_47# VSS 0.01fF
C16884 sky130_fd_sc_hd__dfrtn_1_8/a_1270_413# VSS 0.00fF
C16885 sky130_fd_sc_hd__dfrtn_1_8/a_651_413# VSS 0.02fF
C16886 sky130_fd_sc_hd__dfrtn_1_8/a_448_47# VSS 0.03fF
C16887 sky130_fd_sc_hd__dfrtn_1_8/a_1108_47# VSS 0.21fF
C16888 sky130_fd_sc_hd__dfrtn_1_8/a_1283_21# VSS 0.35fF
C16889 sky130_fd_sc_hd__dfrtn_1_8/a_543_47# VSS 0.18fF
C16890 sky130_fd_sc_hd__dfrtn_1_8/a_761_289# VSS 0.15fF
C16891 sky130_fd_sc_hd__dfrtn_1_8/a_193_47# VSS 0.21fF
C16892 sky130_fd_sc_hd__dfrtn_1_8/a_27_47# VSS 0.49fF
C16893 sky130_fd_sc_hd__nor3_1_3/a_193_297# VSS 0.00fF
C16894 sky130_fd_sc_hd__nor3_1_3/a_109_297# VSS 0.00fF
C16895 sky130_fd_sc_hd__dfrtn_1_7/a_1462_47# VSS 0.00fF
C16896 sky130_fd_sc_hd__dfrtn_1_7/a_1217_47# VSS 0.00fF
C16897 sky130_fd_sc_hd__dfrtn_1_7/a_805_47# VSS 0.00fF
C16898 sky130_fd_sc_hd__dfrtn_1_7/a_639_47# VSS 0.00fF
C16899 sky130_fd_sc_hd__dfrtn_1_7/a_1270_413# VSS 0.00fF
C16900 sky130_fd_sc_hd__dfrtn_1_7/a_651_413# VSS 0.01fF
C16901 sky130_fd_sc_hd__dfrtn_1_7/a_448_47# VSS 0.02fF
C16902 sky130_fd_sc_hd__dfrtn_1_7/a_1108_47# VSS 0.16fF
C16903 sky130_fd_sc_hd__dfrtn_1_7/a_1283_21# VSS 0.31fF
C16904 sky130_fd_sc_hd__dfrtn_1_7/a_543_47# VSS 0.16fF
C16905 sky130_fd_sc_hd__dfrtn_1_7/a_761_289# VSS 0.13fF
C16906 sky130_fd_sc_hd__dfrtn_1_7/a_193_47# VSS 0.28fF
C16907 sky130_fd_sc_hd__dfrtn_1_7/a_27_47# VSS 0.52fF
C16908 sky130_fd_sc_hd__nor3_1_2/a_193_297# VSS 0.00fF
C16909 sky130_fd_sc_hd__nor3_1_2/a_109_297# VSS 0.00fF
C16910 sky130_fd_sc_hd__dfrtn_1_6/a_1462_47# VSS 0.00fF
C16911 sky130_fd_sc_hd__dfrtn_1_6/a_1217_47# VSS 0.00fF
C16912 sky130_fd_sc_hd__dfrtn_1_6/a_805_47# VSS 0.00fF
C16913 sky130_fd_sc_hd__dfrtn_1_6/a_639_47# VSS 0.00fF
C16914 sky130_fd_sc_hd__dfrtn_1_6/a_1270_413# VSS 0.00fF
C16915 sky130_fd_sc_hd__dfrtn_1_6/a_651_413# VSS 0.01fF
C16916 sky130_fd_sc_hd__dfrtn_1_6/a_448_47# VSS 0.02fF
C16917 sky130_fd_sc_hd__dfrtn_1_6/a_1108_47# VSS 0.17fF
C16918 sky130_fd_sc_hd__dfrtn_1_6/a_1283_21# VSS 0.31fF
C16919 sky130_fd_sc_hd__dfrtn_1_6/a_543_47# VSS 0.16fF
C16920 sky130_fd_sc_hd__dfrtn_1_6/a_761_289# VSS 0.13fF
C16921 sky130_fd_sc_hd__dfrtn_1_6/a_193_47# VSS 0.22fF
C16922 sky130_fd_sc_hd__dfrtn_1_6/a_27_47# VSS 0.47fF
C16923 sky130_fd_sc_hd__inv_1_14/A VSS 0.34fF
C16924 sky130_fd_sc_hd__o221ai_1_0/a_213_123# VSS 0.05fF
C16925 sky130_fd_sc_hd__o221ai_1_0/a_109_47# VSS 0.01fF
C16926 sky130_fd_sc_hd__o221ai_1_0/a_493_297# VSS 0.00fF
C16927 sky130_fd_sc_hd__o221ai_1_0/a_295_297# VSS 0.00fF
C16928 sky130_fd_sc_hd__nor3_1_1/a_193_297# VSS 0.00fF
C16929 sky130_fd_sc_hd__nor3_1_1/a_109_297# VSS 0.00fF
C16930 sky130_fd_sc_hd__dfrtn_1_5/a_1462_47# VSS 0.00fF
C16931 sky130_fd_sc_hd__dfrtn_1_5/a_1217_47# VSS 0.00fF
C16932 sky130_fd_sc_hd__dfrtn_1_5/a_805_47# VSS 0.00fF
C16933 sky130_fd_sc_hd__dfrtn_1_5/a_639_47# VSS 0.00fF
C16934 sky130_fd_sc_hd__dfrtn_1_5/a_1270_413# VSS 0.00fF
C16935 sky130_fd_sc_hd__dfrtn_1_5/a_651_413# VSS 0.01fF
C16936 sky130_fd_sc_hd__dfrtn_1_5/a_448_47# VSS 0.02fF
C16937 sky130_fd_sc_hd__dfrtn_1_5/a_1108_47# VSS 0.16fF
C16938 sky130_fd_sc_hd__dfrtn_1_5/a_1283_21# VSS 0.30fF
C16939 sky130_fd_sc_hd__dfrtn_1_5/a_543_47# VSS 0.16fF
C16940 sky130_fd_sc_hd__dfrtn_1_5/a_761_289# VSS 0.13fF
C16941 sky130_fd_sc_hd__dfrtn_1_5/a_193_47# VSS 0.21fF
C16942 sky130_fd_sc_hd__dfrtn_1_5/a_27_47# VSS 0.46fF
C16943 sky130_fd_sc_hd__nor3_1_0/a_193_297# VSS 0.00fF
C16944 sky130_fd_sc_hd__nor3_1_0/a_109_297# VSS 0.00fF
C16945 sky130_fd_sc_hd__dfrtn_1_4/a_1462_47# VSS 0.00fF
C16946 sky130_fd_sc_hd__dfrtn_1_4/a_1217_47# VSS 0.00fF
C16947 sky130_fd_sc_hd__dfrtn_1_4/a_805_47# VSS 0.00fF
C16948 sky130_fd_sc_hd__dfrtn_1_4/a_639_47# VSS 0.00fF
C16949 sky130_fd_sc_hd__dfrtn_1_4/a_1270_413# VSS 0.00fF
C16950 sky130_fd_sc_hd__dfrtn_1_4/a_651_413# VSS 0.01fF
C16951 sky130_fd_sc_hd__dfrtn_1_4/a_448_47# VSS 0.02fF
C16952 sky130_fd_sc_hd__dfrtn_1_4/a_1108_47# VSS 0.17fF
C16953 sky130_fd_sc_hd__dfrtn_1_4/a_1283_21# VSS 0.31fF
C16954 sky130_fd_sc_hd__dfrtn_1_4/a_543_47# VSS 0.16fF
C16955 sky130_fd_sc_hd__dfrtn_1_4/a_761_289# VSS 0.13fF
C16956 sky130_fd_sc_hd__dfrtn_1_4/a_193_47# VSS 0.16fF
C16957 sky130_fd_sc_hd__dfrtn_1_4/a_27_47# VSS 0.44fF
C16958 sky130_fd_sc_hd__dfrtn_1_19/a_1462_47# VSS 0.00fF
C16959 sky130_fd_sc_hd__dfrtn_1_19/a_1217_47# VSS 0.00fF
C16960 sky130_fd_sc_hd__dfrtn_1_19/a_805_47# VSS 0.00fF
C16961 sky130_fd_sc_hd__dfrtn_1_19/a_639_47# VSS 0.00fF
C16962 sky130_fd_sc_hd__dfrtn_1_19/a_1270_413# VSS 0.00fF
C16963 sky130_fd_sc_hd__dfrtn_1_19/a_651_413# VSS 0.01fF
C16964 sky130_fd_sc_hd__dfrtn_1_19/a_448_47# VSS 0.02fF
C16965 sky130_fd_sc_hd__dfrtn_1_19/a_1108_47# VSS 0.15fF
C16966 sky130_fd_sc_hd__dfrtn_1_19/a_1283_21# VSS 0.29fF
C16967 sky130_fd_sc_hd__dfrtn_1_19/a_543_47# VSS 0.15fF
C16968 sky130_fd_sc_hd__dfrtn_1_19/a_761_289# VSS 0.12fF
C16969 sky130_fd_sc_hd__dfrtn_1_19/a_193_47# VSS 0.24fF
C16970 sky130_fd_sc_hd__dfrtn_1_19/a_27_47# VSS 0.44fF
C16971 sky130_fd_sc_hd__nand2_1_2/a_113_47# VSS 0.00fF
C16972 sky130_fd_sc_hd__dfrtn_1_3/a_1462_47# VSS 0.01fF
C16973 sky130_fd_sc_hd__dfrtn_1_3/a_1217_47# VSS 0.00fF
C16974 sky130_fd_sc_hd__dfrtn_1_3/a_805_47# VSS 0.00fF
C16975 sky130_fd_sc_hd__dfrtn_1_3/a_639_47# VSS 0.00fF
C16976 sky130_fd_sc_hd__dfrtn_1_3/a_1270_413# VSS 0.00fF
C16977 sky130_fd_sc_hd__dfrtn_1_3/a_651_413# VSS 0.01fF
C16978 sky130_fd_sc_hd__dfrtn_1_3/a_448_47# VSS 0.02fF
C16979 sky130_fd_sc_hd__dfrtn_1_3/a_1108_47# VSS 0.19fF
C16980 sky130_fd_sc_hd__dfrtn_1_3/a_1283_21# VSS 0.35fF
C16981 sky130_fd_sc_hd__dfrtn_1_3/a_543_47# VSS 0.16fF
C16982 sky130_fd_sc_hd__dfrtn_1_3/a_761_289# VSS 0.13fF
C16983 sky130_fd_sc_hd__dfrtn_1_3/a_193_47# VSS 0.17fF
C16984 sky130_fd_sc_hd__dfrtn_1_3/a_27_47# VSS 0.47fF
C16985 sky130_fd_sc_hd__dfrtn_1_18/a_1462_47# VSS 0.00fF
C16986 sky130_fd_sc_hd__dfrtn_1_18/a_1217_47# VSS 0.00fF
C16987 sky130_fd_sc_hd__dfrtn_1_18/a_805_47# VSS 0.00fF
C16988 sky130_fd_sc_hd__dfrtn_1_18/a_639_47# VSS 0.00fF
C16989 sky130_fd_sc_hd__dfrtn_1_18/a_1270_413# VSS 0.00fF
C16990 sky130_fd_sc_hd__dfrtn_1_18/a_651_413# VSS 0.01fF
C16991 sky130_fd_sc_hd__dfrtn_1_18/a_448_47# VSS 0.01fF
C16992 sky130_fd_sc_hd__dfrtn_1_18/a_1108_47# VSS 0.15fF
C16993 sky130_fd_sc_hd__dfrtn_1_18/a_1283_21# VSS 0.29fF
C16994 sky130_fd_sc_hd__dfrtn_1_18/a_543_47# VSS 0.15fF
C16995 sky130_fd_sc_hd__dfrtn_1_18/a_761_289# VSS 0.12fF
C16996 sky130_fd_sc_hd__dfrtn_1_18/a_193_47# VSS 0.16fF
C16997 sky130_fd_sc_hd__dfrtn_1_18/a_27_47# VSS 0.43fF
C16998 sky130_fd_sc_hd__dfrtn_1_29/a_1462_47# VSS 0.00fF
C16999 sky130_fd_sc_hd__dfrtn_1_29/a_1217_47# VSS 0.00fF
C17000 sky130_fd_sc_hd__dfrtn_1_29/a_805_47# VSS 0.00fF
C17001 sky130_fd_sc_hd__dfrtn_1_29/a_639_47# VSS 0.00fF
C17002 sky130_fd_sc_hd__dfrtn_1_29/a_1270_413# VSS 0.00fF
C17003 sky130_fd_sc_hd__dfrtn_1_29/a_651_413# VSS 0.01fF
C17004 sky130_fd_sc_hd__dfrtn_1_29/a_448_47# VSS 0.02fF
C17005 sky130_fd_sc_hd__dfrtn_1_29/a_1108_47# VSS 0.18fF
C17006 sky130_fd_sc_hd__dfrtn_1_29/a_1283_21# VSS 0.32fF
C17007 sky130_fd_sc_hd__dfrtn_1_29/a_543_47# VSS 0.16fF
C17008 sky130_fd_sc_hd__dfrtn_1_29/a_761_289# VSS 0.13fF
C17009 sky130_fd_sc_hd__dfrtn_1_29/a_193_47# VSS 0.16fF
C17010 sky130_fd_sc_hd__dfrtn_1_29/a_27_47# VSS 0.46fF
C17011 sky130_fd_sc_hd__nand2_1_1/a_113_47# VSS 0.00fF
C17012 sky130_fd_sc_hd__o311a_1_0/a_585_47# VSS 0.00fF
C17013 sky130_fd_sc_hd__o311a_1_0/a_266_47# VSS 0.02fF
C17014 sky130_fd_sc_hd__o311a_1_0/a_368_297# VSS 0.00fF
C17015 sky130_fd_sc_hd__o311a_1_0/a_266_297# VSS 0.00fF
C17016 sky130_fd_sc_hd__o311a_1_0/a_81_21# VSS 0.26fF
C17017 sky130_fd_sc_hd__inv_1_45/Y VSS 0.12fF
C17018 sky130_fd_sc_hd__dfrtn_1_2/a_1462_47# VSS 0.00fF
C17019 sky130_fd_sc_hd__dfrtn_1_2/a_1217_47# VSS 0.00fF
C17020 sky130_fd_sc_hd__dfrtn_1_2/a_805_47# VSS 0.00fF
C17021 sky130_fd_sc_hd__dfrtn_1_2/a_639_47# VSS 0.00fF
C17022 sky130_fd_sc_hd__dfrtn_1_2/a_1270_413# VSS 0.00fF
C17023 sky130_fd_sc_hd__dfrtn_1_2/a_651_413# VSS 0.01fF
C17024 sky130_fd_sc_hd__dfrtn_1_2/a_448_47# VSS 0.02fF
C17025 sky130_fd_sc_hd__dfrtn_1_2/a_1108_47# VSS 0.15fF
C17026 sky130_fd_sc_hd__dfrtn_1_2/a_1283_21# VSS 0.29fF
C17027 sky130_fd_sc_hd__dfrtn_1_2/a_543_47# VSS 0.15fF
C17028 sky130_fd_sc_hd__dfrtn_1_2/a_761_289# VSS 0.12fF
C17029 sky130_fd_sc_hd__dfrtn_1_2/a_193_47# VSS 0.21fF
C17030 sky130_fd_sc_hd__dfrtn_1_2/a_27_47# VSS 0.49fF
C17031 sky130_fd_sc_hd__or2_2_0/a_121_297# VSS 0.00fF
C17032 sky130_fd_sc_hd__or2_2_0/a_39_297# VSS 0.26fF
C17033 sky130_fd_sc_hd__dfrtn_1_17/a_1462_47# VSS 0.00fF
C17034 sky130_fd_sc_hd__dfrtn_1_17/a_1217_47# VSS 0.00fF
C17035 sky130_fd_sc_hd__dfrtn_1_17/a_805_47# VSS 0.00fF
C17036 sky130_fd_sc_hd__dfrtn_1_17/a_639_47# VSS 0.00fF
C17037 sky130_fd_sc_hd__dfrtn_1_17/a_1270_413# VSS 0.00fF
C17038 sky130_fd_sc_hd__dfrtn_1_17/a_651_413# VSS 0.01fF
C17039 sky130_fd_sc_hd__dfrtn_1_17/a_448_47# VSS 0.01fF
C17040 sky130_fd_sc_hd__dfrtn_1_17/a_1108_47# VSS 0.15fF
C17041 sky130_fd_sc_hd__dfrtn_1_17/a_1283_21# VSS 0.29fF
C17042 sky130_fd_sc_hd__dfrtn_1_17/a_543_47# VSS 0.15fF
C17043 sky130_fd_sc_hd__dfrtn_1_17/a_761_289# VSS 0.12fF
C17044 sky130_fd_sc_hd__dfrtn_1_17/a_193_47# VSS 0.23fF
C17045 sky130_fd_sc_hd__dfrtn_1_17/a_27_47# VSS 0.43fF
C17046 sky130_fd_sc_hd__dfrtn_1_28/a_1462_47# VSS 0.00fF
C17047 sky130_fd_sc_hd__dfrtn_1_28/a_1217_47# VSS 0.00fF
C17048 sky130_fd_sc_hd__dfrtn_1_28/a_805_47# VSS 0.00fF
C17049 sky130_fd_sc_hd__dfrtn_1_28/a_639_47# VSS 0.00fF
C17050 sky130_fd_sc_hd__dfrtn_1_28/a_1270_413# VSS 0.00fF
C17051 sky130_fd_sc_hd__dfrtn_1_28/a_651_413# VSS 0.01fF
C17052 sky130_fd_sc_hd__dfrtn_1_28/a_448_47# VSS 0.02fF
C17053 sky130_fd_sc_hd__dfrtn_1_28/a_1108_47# VSS 0.19fF
C17054 sky130_fd_sc_hd__dfrtn_1_28/a_1283_21# VSS 0.33fF
C17055 sky130_fd_sc_hd__dfrtn_1_28/a_543_47# VSS 0.17fF
C17056 sky130_fd_sc_hd__dfrtn_1_28/a_761_289# VSS 0.14fF
C17057 sky130_fd_sc_hd__dfrtn_1_28/a_193_47# VSS 0.19fF
C17058 sky130_fd_sc_hd__dfrtn_1_28/a_27_47# VSS 0.47fF
C17059 sky130_fd_sc_hd__dfrtn_1_39/a_1462_47# VSS 0.00fF
C17060 sky130_fd_sc_hd__dfrtn_1_39/a_1217_47# VSS 0.00fF
C17061 sky130_fd_sc_hd__dfrtn_1_39/a_805_47# VSS 0.00fF
C17062 sky130_fd_sc_hd__dfrtn_1_39/a_639_47# VSS 0.00fF
C17063 sky130_fd_sc_hd__dfrtn_1_39/a_1270_413# VSS 0.00fF
C17064 sky130_fd_sc_hd__dfrtn_1_39/a_651_413# VSS 0.01fF
C17065 sky130_fd_sc_hd__dfrtn_1_39/a_448_47# VSS 0.01fF
C17066 sky130_fd_sc_hd__dfrtn_1_39/a_1108_47# VSS 0.15fF
C17067 sky130_fd_sc_hd__dfrtn_1_39/a_1283_21# VSS 0.29fF
C17068 sky130_fd_sc_hd__dfrtn_1_39/a_543_47# VSS 0.15fF
C17069 sky130_fd_sc_hd__dfrtn_1_39/a_761_289# VSS 0.12fF
C17070 sky130_fd_sc_hd__dfrtn_1_39/a_193_47# VSS 0.25fF
C17071 sky130_fd_sc_hd__dfrtn_1_39/a_27_47# VSS 0.43fF
C17072 DOUT[9] VSS 8.95fF
C17073 sky130_fd_sc_hd__nand2_1_0/a_113_47# VSS 0.00fF
C17074 sky130_fd_sc_hd__mux4_2_0/a_1281_47# VSS 0.00fF
C17075 sky130_fd_sc_hd__mux4_2_0/a_1064_47# VSS 0.00fF
C17076 sky130_fd_sc_hd__mux4_2_0/a_397_47# VSS 0.00fF
C17077 sky130_fd_sc_hd__mux4_2_0/a_1279_413# VSS -0.00fF
C17078 sky130_fd_sc_hd__mux4_2_0/a_1060_369# VSS -0.00fF
C17079 sky130_fd_sc_hd__mux4_2_0/a_872_316# VSS 0.04fF
C17080 sky130_fd_sc_hd__mux4_2_0/a_193_47# VSS 0.00fF
C17081 sky130_fd_sc_hd__mux4_2_0/a_600_345# VSS 0.11fF
C17082 sky130_fd_sc_hd__mux4_2_0/a_788_316# VSS 0.23fF
C17083 sky130_fd_sc_hd__mux4_2_0/a_372_413# VSS 0.00fF
C17084 sky130_fd_sc_hd__mux4_2_0/a_288_47# VSS 0.03fF
C17085 sky130_fd_sc_hd__mux4_2_0/a_193_369# VSS 0.00fF
C17086 sky130_fd_sc_hd__mux4_2_0/a_27_47# VSS 0.29fF
C17087 sky130_fd_sc_hd__dfrtn_1_1/a_1462_47# VSS 0.00fF
C17088 sky130_fd_sc_hd__dfrtn_1_1/a_1217_47# VSS 0.00fF
C17089 sky130_fd_sc_hd__dfrtn_1_1/a_805_47# VSS 0.00fF
C17090 sky130_fd_sc_hd__dfrtn_1_1/a_639_47# VSS 0.00fF
C17091 sky130_fd_sc_hd__dfrtn_1_1/a_1270_413# VSS 0.00fF
C17092 sky130_fd_sc_hd__dfrtn_1_1/a_651_413# VSS 0.01fF
C17093 sky130_fd_sc_hd__dfrtn_1_1/a_448_47# VSS 0.02fF
C17094 sky130_fd_sc_hd__dfrtn_1_1/a_1108_47# VSS 0.17fF
C17095 sky130_fd_sc_hd__dfrtn_1_1/a_1283_21# VSS 0.31fF
C17096 sky130_fd_sc_hd__dfrtn_1_1/a_543_47# VSS 0.16fF
C17097 sky130_fd_sc_hd__dfrtn_1_1/a_761_289# VSS 0.12fF
C17098 sky130_fd_sc_hd__dfrtn_1_1/a_193_47# VSS 0.18fF
C17099 sky130_fd_sc_hd__dfrtn_1_1/a_27_47# VSS 0.43fF
C17100 sky130_fd_sc_hd__dfrtn_1_16/a_1462_47# VSS 0.00fF
C17101 sky130_fd_sc_hd__dfrtn_1_16/a_1217_47# VSS 0.00fF
C17102 sky130_fd_sc_hd__dfrtn_1_16/a_805_47# VSS 0.00fF
C17103 sky130_fd_sc_hd__dfrtn_1_16/a_639_47# VSS 0.00fF
C17104 sky130_fd_sc_hd__dfrtn_1_16/a_1270_413# VSS 0.00fF
C17105 sky130_fd_sc_hd__dfrtn_1_16/a_651_413# VSS 0.01fF
C17106 sky130_fd_sc_hd__dfrtn_1_16/a_448_47# VSS 0.02fF
C17107 sky130_fd_sc_hd__dfrtn_1_16/a_1108_47# VSS 0.15fF
C17108 sky130_fd_sc_hd__dfrtn_1_16/a_1283_21# VSS 0.29fF
C17109 sky130_fd_sc_hd__dfrtn_1_16/a_543_47# VSS 0.15fF
C17110 sky130_fd_sc_hd__dfrtn_1_16/a_761_289# VSS 0.12fF
C17111 sky130_fd_sc_hd__dfrtn_1_16/a_193_47# VSS 0.15fF
C17112 sky130_fd_sc_hd__dfrtn_1_16/a_27_47# VSS 0.43fF
C17113 sky130_fd_sc_hd__dfrtn_1_27/a_1462_47# VSS 0.00fF
C17114 sky130_fd_sc_hd__dfrtn_1_27/a_1217_47# VSS 0.00fF
C17115 sky130_fd_sc_hd__dfrtn_1_27/a_805_47# VSS 0.00fF
C17116 sky130_fd_sc_hd__dfrtn_1_27/a_639_47# VSS 0.00fF
C17117 sky130_fd_sc_hd__dfrtn_1_27/a_1270_413# VSS 0.00fF
C17118 sky130_fd_sc_hd__dfrtn_1_27/a_651_413# VSS 0.00fF
C17119 sky130_fd_sc_hd__dfrtn_1_27/a_448_47# VSS 0.01fF
C17120 sky130_fd_sc_hd__dfrtn_1_27/a_1108_47# VSS 0.15fF
C17121 sky130_fd_sc_hd__dfrtn_1_27/a_1283_21# VSS 0.29fF
C17122 sky130_fd_sc_hd__dfrtn_1_27/a_543_47# VSS 0.14fF
C17123 sky130_fd_sc_hd__dfrtn_1_27/a_761_289# VSS 0.11fF
C17124 sky130_fd_sc_hd__dfrtn_1_27/a_193_47# VSS 0.14fF
C17125 sky130_fd_sc_hd__dfrtn_1_27/a_27_47# VSS 0.42fF
C17126 sky130_fd_sc_hd__dfrtn_1_38/a_1462_47# VSS 0.00fF
C17127 sky130_fd_sc_hd__dfrtn_1_38/a_1217_47# VSS 0.00fF
C17128 sky130_fd_sc_hd__dfrtn_1_38/a_805_47# VSS 0.00fF
C17129 sky130_fd_sc_hd__dfrtn_1_38/a_639_47# VSS 0.00fF
C17130 sky130_fd_sc_hd__dfrtn_1_38/a_1270_413# VSS 0.00fF
C17131 sky130_fd_sc_hd__dfrtn_1_38/a_651_413# VSS 0.01fF
C17132 sky130_fd_sc_hd__dfrtn_1_38/a_448_47# VSS 0.01fF
C17133 sky130_fd_sc_hd__dfrtn_1_38/a_1108_47# VSS 0.15fF
C17134 sky130_fd_sc_hd__dfrtn_1_38/a_1283_21# VSS 0.29fF
C17135 sky130_fd_sc_hd__dfrtn_1_38/a_543_47# VSS 0.15fF
C17136 sky130_fd_sc_hd__dfrtn_1_38/a_761_289# VSS 0.12fF
C17137 sky130_fd_sc_hd__dfrtn_1_38/a_193_47# VSS 0.22fF
C17138 sky130_fd_sc_hd__dfrtn_1_38/a_27_47# VSS 0.45fF
C17139 sky130_fd_sc_hd__dfrtn_1_0/a_1462_47# VSS 0.00fF
C17140 sky130_fd_sc_hd__dfrtn_1_0/a_1217_47# VSS 0.00fF
C17141 sky130_fd_sc_hd__dfrtn_1_0/a_805_47# VSS 0.00fF
C17142 sky130_fd_sc_hd__dfrtn_1_0/a_639_47# VSS 0.00fF
C17143 sky130_fd_sc_hd__dfrtn_1_0/a_1270_413# VSS 0.00fF
C17144 sky130_fd_sc_hd__dfrtn_1_0/a_651_413# VSS 0.01fF
C17145 sky130_fd_sc_hd__dfrtn_1_0/a_448_47# VSS 0.02fF
C17146 sky130_fd_sc_hd__dfrtn_1_0/a_1108_47# VSS 0.16fF
C17147 sky130_fd_sc_hd__dfrtn_1_0/a_1283_21# VSS 0.30fF
C17148 sky130_fd_sc_hd__dfrtn_1_0/a_543_47# VSS 0.16fF
C17149 sky130_fd_sc_hd__dfrtn_1_0/a_761_289# VSS 0.13fF
C17150 sky130_fd_sc_hd__dfrtn_1_0/a_193_47# VSS 0.21fF
C17151 sky130_fd_sc_hd__dfrtn_1_0/a_27_47# VSS 0.45fF
C17152 sky130_fd_sc_hd__dfrtn_1_15/a_1462_47# VSS 0.00fF
C17153 sky130_fd_sc_hd__dfrtn_1_15/a_1217_47# VSS 0.00fF
C17154 sky130_fd_sc_hd__dfrtn_1_15/a_805_47# VSS 0.00fF
C17155 sky130_fd_sc_hd__dfrtn_1_15/a_639_47# VSS 0.00fF
C17156 sky130_fd_sc_hd__dfrtn_1_15/a_1270_413# VSS 0.00fF
C17157 sky130_fd_sc_hd__dfrtn_1_15/a_651_413# VSS 0.01fF
C17158 sky130_fd_sc_hd__dfrtn_1_15/a_448_47# VSS 0.02fF
C17159 sky130_fd_sc_hd__dfrtn_1_15/a_1108_47# VSS 0.16fF
C17160 sky130_fd_sc_hd__dfrtn_1_15/a_1283_21# VSS 0.30fF
C17161 sky130_fd_sc_hd__dfrtn_1_15/a_543_47# VSS 0.16fF
C17162 sky130_fd_sc_hd__dfrtn_1_15/a_761_289# VSS 0.13fF
C17163 sky130_fd_sc_hd__dfrtn_1_15/a_193_47# VSS 0.19fF
C17164 sky130_fd_sc_hd__dfrtn_1_15/a_27_47# VSS 0.47fF
C17165 sky130_fd_sc_hd__dfrtn_1_26/a_1462_47# VSS 0.00fF
C17166 sky130_fd_sc_hd__dfrtn_1_26/a_1217_47# VSS 0.00fF
C17167 sky130_fd_sc_hd__dfrtn_1_26/a_805_47# VSS 0.00fF
C17168 sky130_fd_sc_hd__dfrtn_1_26/a_639_47# VSS 0.00fF
C17169 sky130_fd_sc_hd__dfrtn_1_26/a_1270_413# VSS 0.00fF
C17170 sky130_fd_sc_hd__dfrtn_1_26/a_651_413# VSS 0.01fF
C17171 sky130_fd_sc_hd__dfrtn_1_26/a_448_47# VSS 0.01fF
C17172 sky130_fd_sc_hd__dfrtn_1_26/a_1108_47# VSS 0.15fF
C17173 sky130_fd_sc_hd__dfrtn_1_26/a_1283_21# VSS 0.29fF
C17174 sky130_fd_sc_hd__dfrtn_1_26/a_543_47# VSS 0.15fF
C17175 sky130_fd_sc_hd__dfrtn_1_26/a_761_289# VSS 0.12fF
C17176 sky130_fd_sc_hd__dfrtn_1_26/a_193_47# VSS 0.14fF
C17177 sky130_fd_sc_hd__dfrtn_1_26/a_27_47# VSS 0.42fF
C17178 sky130_fd_sc_hd__dfrtn_1_37/a_1462_47# VSS 0.00fF
C17179 sky130_fd_sc_hd__dfrtn_1_37/a_1217_47# VSS 0.00fF
C17180 sky130_fd_sc_hd__dfrtn_1_37/a_805_47# VSS 0.00fF
C17181 sky130_fd_sc_hd__dfrtn_1_37/a_639_47# VSS 0.00fF
C17182 sky130_fd_sc_hd__dfrtn_1_37/a_1270_413# VSS 0.00fF
C17183 sky130_fd_sc_hd__dfrtn_1_37/a_651_413# VSS 0.01fF
C17184 sky130_fd_sc_hd__dfrtn_1_37/a_448_47# VSS 0.01fF
C17185 sky130_fd_sc_hd__dfrtn_1_37/a_1108_47# VSS 0.15fF
C17186 sky130_fd_sc_hd__dfrtn_1_37/a_1283_21# VSS 0.28fF
C17187 sky130_fd_sc_hd__dfrtn_1_37/a_543_47# VSS 0.15fF
C17188 sky130_fd_sc_hd__dfrtn_1_37/a_761_289# VSS 0.12fF
C17189 sky130_fd_sc_hd__dfrtn_1_37/a_193_47# VSS 0.14fF
C17190 sky130_fd_sc_hd__dfrtn_1_37/a_27_47# VSS 0.42fF
C17191 sky130_fd_sc_hd__conb_1_0/LO VSS 0.23fF
C17192 sky130_fd_sc_hd__dfrtn_1_36/a_1462_47# VSS 0.00fF
C17193 sky130_fd_sc_hd__dfrtn_1_36/a_1217_47# VSS 0.00fF
C17194 sky130_fd_sc_hd__dfrtn_1_36/a_805_47# VSS 0.00fF
C17195 sky130_fd_sc_hd__dfrtn_1_36/a_639_47# VSS 0.00fF
C17196 sky130_fd_sc_hd__dfrtn_1_36/a_1270_413# VSS 0.00fF
C17197 sky130_fd_sc_hd__dfrtn_1_36/a_651_413# VSS 0.01fF
C17198 sky130_fd_sc_hd__dfrtn_1_36/a_448_47# VSS 0.02fF
C17199 sky130_fd_sc_hd__dfrtn_1_36/a_1108_47# VSS 0.18fF
C17200 sky130_fd_sc_hd__dfrtn_1_36/a_1283_21# VSS 0.29fF
C17201 sky130_fd_sc_hd__dfrtn_1_36/a_543_47# VSS 0.17fF
C17202 sky130_fd_sc_hd__dfrtn_1_36/a_761_289# VSS 0.14fF
C17203 sky130_fd_sc_hd__dfrtn_1_36/a_193_47# VSS 0.20fF
C17204 sky130_fd_sc_hd__dfrtn_1_36/a_27_47# VSS 0.49fF
C17205 sky130_fd_sc_hd__dfrtn_1_14/a_1462_47# VSS 0.00fF
C17206 sky130_fd_sc_hd__dfrtn_1_14/a_1217_47# VSS 0.00fF
C17207 sky130_fd_sc_hd__dfrtn_1_14/a_805_47# VSS 0.00fF
C17208 sky130_fd_sc_hd__dfrtn_1_14/a_639_47# VSS 0.00fF
C17209 sky130_fd_sc_hd__dfrtn_1_14/a_1270_413# VSS 0.00fF
C17210 sky130_fd_sc_hd__dfrtn_1_14/a_651_413# VSS 0.01fF
C17211 sky130_fd_sc_hd__dfrtn_1_14/a_448_47# VSS 0.01fF
C17212 sky130_fd_sc_hd__dfrtn_1_14/a_1108_47# VSS 0.15fF
C17213 sky130_fd_sc_hd__dfrtn_1_14/a_1283_21# VSS 0.28fF
C17214 sky130_fd_sc_hd__dfrtn_1_14/a_543_47# VSS 0.15fF
C17215 sky130_fd_sc_hd__dfrtn_1_14/a_761_289# VSS 0.12fF
C17216 sky130_fd_sc_hd__dfrtn_1_14/a_193_47# VSS 0.16fF
C17217 sky130_fd_sc_hd__dfrtn_1_14/a_27_47# VSS 0.50fF
C17218 sky130_fd_sc_hd__dfrtn_1_25/a_1462_47# VSS 0.00fF
C17219 sky130_fd_sc_hd__dfrtn_1_25/a_1217_47# VSS 0.00fF
C17220 sky130_fd_sc_hd__dfrtn_1_25/a_805_47# VSS 0.00fF
C17221 sky130_fd_sc_hd__dfrtn_1_25/a_639_47# VSS 0.00fF
C17222 sky130_fd_sc_hd__dfrtn_1_25/a_1270_413# VSS 0.00fF
C17223 sky130_fd_sc_hd__dfrtn_1_25/a_651_413# VSS 0.01fF
C17224 sky130_fd_sc_hd__dfrtn_1_25/a_448_47# VSS 0.01fF
C17225 sky130_fd_sc_hd__dfrtn_1_25/a_1108_47# VSS 0.16fF
C17226 sky130_fd_sc_hd__dfrtn_1_25/a_1283_21# VSS 0.30fF
C17227 sky130_fd_sc_hd__dfrtn_1_25/a_543_47# VSS 0.15fF
C17228 sky130_fd_sc_hd__dfrtn_1_25/a_761_289# VSS 0.12fF
C17229 sky130_fd_sc_hd__dfrtn_1_25/a_193_47# VSS 0.26fF
C17230 sky130_fd_sc_hd__dfrtn_1_25/a_27_47# VSS 0.45fF
C17231 sky130_fd_sc_hd__inv_1_21/Y VSS 0.25fF
C17232 sky130_fd_sc_hd__inv_1_45/A VSS 0.38fF
C17233 sky130_fd_sc_hd__dfrtn_1_13/a_1462_47# VSS 0.00fF
C17234 sky130_fd_sc_hd__dfrtn_1_13/a_1217_47# VSS 0.00fF
C17235 sky130_fd_sc_hd__dfrtn_1_13/a_805_47# VSS 0.00fF
C17236 sky130_fd_sc_hd__dfrtn_1_13/a_639_47# VSS 0.01fF
C17237 sky130_fd_sc_hd__dfrtn_1_13/a_1270_413# VSS 0.00fF
C17238 sky130_fd_sc_hd__dfrtn_1_13/a_651_413# VSS 0.01fF
C17239 sky130_fd_sc_hd__dfrtn_1_13/a_448_47# VSS 0.02fF
C17240 sky130_fd_sc_hd__dfrtn_1_13/a_1108_47# VSS 0.18fF
C17241 sky130_fd_sc_hd__dfrtn_1_13/a_1283_21# VSS 0.35fF
C17242 sky130_fd_sc_hd__dfrtn_1_13/a_543_47# VSS 0.18fF
C17243 sky130_fd_sc_hd__dfrtn_1_13/a_761_289# VSS 0.14fF
C17244 sky130_fd_sc_hd__dfrtn_1_13/a_193_47# VSS 0.29fF
C17245 sky130_fd_sc_hd__dfrtn_1_13/a_27_47# VSS 0.52fF
C17246 sky130_fd_sc_hd__dfrtn_1_35/a_1462_47# VSS 0.00fF
C17247 sky130_fd_sc_hd__dfrtn_1_35/a_1217_47# VSS 0.00fF
C17248 sky130_fd_sc_hd__dfrtn_1_35/a_805_47# VSS 0.00fF
C17249 sky130_fd_sc_hd__dfrtn_1_35/a_639_47# VSS 0.01fF
C17250 sky130_fd_sc_hd__dfrtn_1_35/a_1270_413# VSS 0.00fF
C17251 sky130_fd_sc_hd__dfrtn_1_35/a_651_413# VSS 0.01fF
C17252 sky130_fd_sc_hd__dfrtn_1_35/a_448_47# VSS 0.04fF
C17253 sky130_fd_sc_hd__dfrtn_1_35/a_1108_47# VSS 0.16fF
C17254 sky130_fd_sc_hd__dfrtn_1_35/a_1283_21# VSS 0.30fF
C17255 sky130_fd_sc_hd__dfrtn_1_35/a_543_47# VSS 0.19fF
C17256 sky130_fd_sc_hd__dfrtn_1_35/a_761_289# VSS 0.13fF
C17257 sky130_fd_sc_hd__dfrtn_1_35/a_193_47# VSS 0.31fF
C17258 sky130_fd_sc_hd__dfrtn_1_35/a_27_47# VSS 0.54fF
C17259 sky130_fd_sc_hd__dfrtn_1_24/a_1462_47# VSS 0.00fF
C17260 sky130_fd_sc_hd__dfrtn_1_24/a_1217_47# VSS 0.00fF
C17261 sky130_fd_sc_hd__dfrtn_1_24/a_805_47# VSS 0.00fF
C17262 sky130_fd_sc_hd__dfrtn_1_24/a_639_47# VSS 0.00fF
C17263 sky130_fd_sc_hd__dfrtn_1_24/a_1270_413# VSS 0.00fF
C17264 sky130_fd_sc_hd__dfrtn_1_24/a_651_413# VSS 0.01fF
C17265 sky130_fd_sc_hd__dfrtn_1_24/a_448_47# VSS 0.02fF
C17266 sky130_fd_sc_hd__dfrtn_1_24/a_1108_47# VSS 0.16fF
C17267 sky130_fd_sc_hd__dfrtn_1_24/a_1283_21# VSS 0.29fF
C17268 sky130_fd_sc_hd__dfrtn_1_24/a_543_47# VSS 0.16fF
C17269 sky130_fd_sc_hd__dfrtn_1_24/a_761_289# VSS 0.13fF
C17270 sky130_fd_sc_hd__dfrtn_1_24/a_193_47# VSS 0.19fF
C17271 sky130_fd_sc_hd__dfrtn_1_24/a_27_47# VSS 0.51fF
C17272 sky130_fd_sc_hd__o211a_1_1/a_510_47# VSS 0.00fF
C17273 sky130_fd_sc_hd__o211a_1_1/a_215_47# VSS 0.02fF
C17274 sky130_fd_sc_hd__o211a_1_1/a_297_297# VSS 0.00fF
C17275 sky130_fd_sc_hd__o211a_1_1/a_79_21# VSS 0.28fF
C17276 sky130_fd_sc_hd__dfrtn_1_23/a_1462_47# VSS 0.00fF
C17277 sky130_fd_sc_hd__dfrtn_1_23/a_1217_47# VSS 0.00fF
C17278 sky130_fd_sc_hd__dfrtn_1_23/a_805_47# VSS 0.00fF
C17279 sky130_fd_sc_hd__dfrtn_1_23/a_639_47# VSS 0.00fF
C17280 sky130_fd_sc_hd__dfrtn_1_23/a_1270_413# VSS 0.00fF
C17281 sky130_fd_sc_hd__dfrtn_1_23/a_651_413# VSS 0.01fF
C17282 sky130_fd_sc_hd__dfrtn_1_23/a_448_47# VSS 0.01fF
C17283 sky130_fd_sc_hd__dfrtn_1_23/a_1108_47# VSS 0.14fF
C17284 sky130_fd_sc_hd__dfrtn_1_23/a_1283_21# VSS 0.28fF
C17285 sky130_fd_sc_hd__dfrtn_1_23/a_543_47# VSS 0.15fF
C17286 sky130_fd_sc_hd__dfrtn_1_23/a_761_289# VSS 0.11fF
C17287 sky130_fd_sc_hd__dfrtn_1_23/a_193_47# VSS 0.14fF
C17288 sky130_fd_sc_hd__dfrtn_1_23/a_27_47# VSS 0.45fF
C17289 sky130_fd_sc_hd__dfrtn_1_12/a_1462_47# VSS 0.00fF
C17290 sky130_fd_sc_hd__dfrtn_1_12/a_1217_47# VSS 0.00fF
C17291 sky130_fd_sc_hd__dfrtn_1_12/a_805_47# VSS 0.00fF
C17292 sky130_fd_sc_hd__dfrtn_1_12/a_639_47# VSS 0.00fF
C17293 sky130_fd_sc_hd__dfrtn_1_12/a_1270_413# VSS 0.00fF
C17294 sky130_fd_sc_hd__dfrtn_1_12/a_651_413# VSS 0.01fF
C17295 sky130_fd_sc_hd__dfrtn_1_12/a_448_47# VSS 0.02fF
C17296 sky130_fd_sc_hd__dfrtn_1_12/a_1108_47# VSS 0.17fF
C17297 sky130_fd_sc_hd__dfrtn_1_12/a_1283_21# VSS 0.31fF
C17298 sky130_fd_sc_hd__dfrtn_1_12/a_543_47# VSS 0.17fF
C17299 sky130_fd_sc_hd__dfrtn_1_12/a_761_289# VSS 0.13fF
C17300 sky130_fd_sc_hd__dfrtn_1_12/a_193_47# VSS 0.17fF
C17301 sky130_fd_sc_hd__dfrtn_1_12/a_27_47# VSS 0.47fF
C17302 sky130_fd_sc_hd__dfrtn_1_34/a_1462_47# VSS 0.00fF
C17303 sky130_fd_sc_hd__dfrtn_1_34/a_1217_47# VSS 0.00fF
C17304 sky130_fd_sc_hd__dfrtn_1_34/a_805_47# VSS 0.00fF
C17305 sky130_fd_sc_hd__dfrtn_1_34/a_639_47# VSS 0.00fF
C17306 sky130_fd_sc_hd__dfrtn_1_34/a_1270_413# VSS 0.00fF
C17307 sky130_fd_sc_hd__dfrtn_1_34/a_651_413# VSS 0.01fF
C17308 sky130_fd_sc_hd__dfrtn_1_34/a_448_47# VSS 0.01fF
C17309 sky130_fd_sc_hd__dfrtn_1_34/a_1108_47# VSS 0.15fF
C17310 sky130_fd_sc_hd__dfrtn_1_34/a_1283_21# VSS 0.28fF
C17311 sky130_fd_sc_hd__dfrtn_1_34/a_543_47# VSS 0.15fF
C17312 sky130_fd_sc_hd__dfrtn_1_34/a_761_289# VSS 0.12fF
C17313 sky130_fd_sc_hd__dfrtn_1_34/a_193_47# VSS 0.21fF
C17314 sky130_fd_sc_hd__dfrtn_1_34/a_27_47# VSS 0.46fF
C17315 sky130_fd_sc_hd__inv_1_46/Y VSS 0.10fF
C17316 sky130_fd_sc_hd__o211a_1_0/a_510_47# VSS 0.00fF
C17317 sky130_fd_sc_hd__o211a_1_0/a_215_47# VSS 0.02fF
C17318 sky130_fd_sc_hd__o211a_1_0/a_297_297# VSS 0.00fF
C17319 sky130_fd_sc_hd__o211a_1_0/a_79_21# VSS 0.27fF
C17320 sky130_fd_sc_hd__dfrtn_1_22/a_1462_47# VSS 0.00fF
C17321 sky130_fd_sc_hd__dfrtn_1_22/a_1217_47# VSS 0.00fF
C17322 sky130_fd_sc_hd__dfrtn_1_22/a_805_47# VSS 0.00fF
C17323 sky130_fd_sc_hd__dfrtn_1_22/a_639_47# VSS 0.00fF
C17324 sky130_fd_sc_hd__dfrtn_1_22/a_1270_413# VSS 0.00fF
C17325 sky130_fd_sc_hd__dfrtn_1_22/a_651_413# VSS 0.01fF
C17326 sky130_fd_sc_hd__dfrtn_1_22/a_448_47# VSS 0.01fF
C17327 sky130_fd_sc_hd__dfrtn_1_22/a_1108_47# VSS 0.16fF
C17328 sky130_fd_sc_hd__dfrtn_1_22/a_1283_21# VSS 0.29fF
C17329 sky130_fd_sc_hd__dfrtn_1_22/a_543_47# VSS 0.15fF
C17330 sky130_fd_sc_hd__dfrtn_1_22/a_761_289# VSS 0.12fF
C17331 sky130_fd_sc_hd__dfrtn_1_22/a_193_47# VSS 0.27fF
C17332 sky130_fd_sc_hd__dfrtn_1_22/a_27_47# VSS 0.44fF
C17333 sky130_fd_sc_hd__dfrtn_1_11/a_1462_47# VSS 0.00fF
C17334 sky130_fd_sc_hd__dfrtn_1_11/a_1217_47# VSS 0.00fF
C17335 sky130_fd_sc_hd__dfrtn_1_11/a_805_47# VSS 0.00fF
C17336 sky130_fd_sc_hd__dfrtn_1_11/a_639_47# VSS 0.00fF
C17337 sky130_fd_sc_hd__dfrtn_1_11/a_1270_413# VSS 0.00fF
C17338 sky130_fd_sc_hd__dfrtn_1_11/a_651_413# VSS 0.01fF
C17339 sky130_fd_sc_hd__dfrtn_1_11/a_448_47# VSS 0.02fF
C17340 sky130_fd_sc_hd__dfrtn_1_11/a_1108_47# VSS 0.15fF
C17341 sky130_fd_sc_hd__dfrtn_1_11/a_1283_21# VSS 0.29fF
C17342 sky130_fd_sc_hd__dfrtn_1_11/a_543_47# VSS 0.15fF
C17343 sky130_fd_sc_hd__dfrtn_1_11/a_761_289# VSS 0.12fF
C17344 sky130_fd_sc_hd__dfrtn_1_11/a_193_47# VSS 0.18fF
C17345 sky130_fd_sc_hd__dfrtn_1_11/a_27_47# VSS 0.45fF
C17346 sky130_fd_sc_hd__dfrtn_1_33/a_1462_47# VSS 0.00fF
C17347 sky130_fd_sc_hd__dfrtn_1_33/a_1217_47# VSS 0.00fF
C17348 sky130_fd_sc_hd__dfrtn_1_33/a_805_47# VSS 0.00fF
C17349 sky130_fd_sc_hd__dfrtn_1_33/a_639_47# VSS 0.00fF
C17350 sky130_fd_sc_hd__dfrtn_1_33/a_1270_413# VSS 0.00fF
C17351 sky130_fd_sc_hd__dfrtn_1_33/a_651_413# VSS 0.01fF
C17352 sky130_fd_sc_hd__dfrtn_1_33/a_448_47# VSS 0.02fF
C17353 sky130_fd_sc_hd__dfrtn_1_33/a_1108_47# VSS 0.16fF
C17354 sky130_fd_sc_hd__dfrtn_1_33/a_1283_21# VSS 0.30fF
C17355 sky130_fd_sc_hd__dfrtn_1_33/a_543_47# VSS 0.16fF
C17356 sky130_fd_sc_hd__dfrtn_1_33/a_761_289# VSS 0.13fF
C17357 sky130_fd_sc_hd__dfrtn_1_33/a_193_47# VSS 0.26fF
C17358 sky130_fd_sc_hd__dfrtn_1_33/a_27_47# VSS 0.44fF
C17359 sky130_fd_sc_hd__inv_1_54/A VSS 0.79fF
C17360 sky130_fd_sc_hd__inv_1_47/Y VSS 0.15fF
C17361 sky130_fd_sc_hd__dfrtn_1_32/a_1462_47# VSS 0.00fF
C17362 sky130_fd_sc_hd__dfrtn_1_32/a_1217_47# VSS 0.00fF
C17363 sky130_fd_sc_hd__dfrtn_1_32/a_805_47# VSS 0.00fF
C17364 sky130_fd_sc_hd__dfrtn_1_32/a_639_47# VSS 0.00fF
C17365 sky130_fd_sc_hd__dfrtn_1_32/a_1270_413# VSS 0.00fF
C17366 sky130_fd_sc_hd__dfrtn_1_32/a_651_413# VSS 0.01fF
C17367 sky130_fd_sc_hd__dfrtn_1_32/a_448_47# VSS 0.01fF
C17368 sky130_fd_sc_hd__dfrtn_1_32/a_1108_47# VSS 0.15fF
C17369 sky130_fd_sc_hd__dfrtn_1_32/a_1283_21# VSS 0.32fF
C17370 sky130_fd_sc_hd__dfrtn_1_32/a_543_47# VSS 0.15fF
C17371 sky130_fd_sc_hd__dfrtn_1_32/a_761_289# VSS 0.12fF
C17372 sky130_fd_sc_hd__dfrtn_1_32/a_193_47# VSS 0.17fF
C17373 sky130_fd_sc_hd__dfrtn_1_32/a_27_47# VSS 0.43fF
C17374 sky130_fd_sc_hd__dfrtn_1_10/a_1462_47# VSS 0.00fF
C17375 sky130_fd_sc_hd__dfrtn_1_10/a_1217_47# VSS 0.00fF
C17376 sky130_fd_sc_hd__dfrtn_1_10/a_805_47# VSS 0.00fF
C17377 sky130_fd_sc_hd__dfrtn_1_10/a_639_47# VSS 0.00fF
C17378 sky130_fd_sc_hd__dfrtn_1_10/a_1270_413# VSS 0.00fF
C17379 sky130_fd_sc_hd__dfrtn_1_10/a_651_413# VSS 0.01fF
C17380 sky130_fd_sc_hd__dfrtn_1_10/a_448_47# VSS 0.02fF
C17381 sky130_fd_sc_hd__dfrtn_1_10/a_1108_47# VSS 0.19fF
C17382 sky130_fd_sc_hd__dfrtn_1_10/a_1283_21# VSS 0.34fF
C17383 sky130_fd_sc_hd__dfrtn_1_10/a_543_47# VSS 0.17fF
C17384 sky130_fd_sc_hd__dfrtn_1_10/a_761_289# VSS 0.14fF
C17385 sky130_fd_sc_hd__dfrtn_1_10/a_193_47# VSS 0.26fF
C17386 sky130_fd_sc_hd__dfrtn_1_10/a_27_47# VSS 0.46fF
C17387 sky130_fd_sc_hd__dfrtn_1_21/a_1462_47# VSS 0.00fF
C17388 sky130_fd_sc_hd__dfrtn_1_21/a_1217_47# VSS 0.00fF
C17389 sky130_fd_sc_hd__dfrtn_1_21/a_805_47# VSS 0.00fF
C17390 sky130_fd_sc_hd__dfrtn_1_21/a_639_47# VSS 0.00fF
C17391 sky130_fd_sc_hd__dfrtn_1_21/a_1270_413# VSS 0.00fF
C17392 sky130_fd_sc_hd__dfrtn_1_21/a_651_413# VSS 0.01fF
C17393 sky130_fd_sc_hd__dfrtn_1_21/a_448_47# VSS 0.01fF
C17394 sky130_fd_sc_hd__dfrtn_1_21/a_1108_47# VSS 0.15fF
C17395 sky130_fd_sc_hd__dfrtn_1_21/a_1283_21# VSS 0.29fF
C17396 sky130_fd_sc_hd__dfrtn_1_21/a_543_47# VSS 0.15fF
C17397 sky130_fd_sc_hd__dfrtn_1_21/a_761_289# VSS 0.12fF
C17398 sky130_fd_sc_hd__dfrtn_1_21/a_193_47# VSS 0.14fF
C17399 sky130_fd_sc_hd__dfrtn_1_21/a_27_47# VSS 0.45fF
C17400 SLC_0/a_1235_416# VSS 0.00fF
C17401 SLC_0/a_919_243# VSS 0.28fF
C17402 SLC_0/a_264_22# VSS 0.33fF
C17403 SLC_0/a_438_293# VSS 0.15fF
C17404 sky130_fd_sc_hd__inv_1_31/A VSS 2.51fF
C17405 sky130_fd_sc_hd__dfrtn_1_42/a_1462_47# VSS 0.00fF
C17406 sky130_fd_sc_hd__dfrtn_1_42/a_1217_47# VSS 0.00fF
C17407 sky130_fd_sc_hd__dfrtn_1_42/a_805_47# VSS 0.00fF
C17408 sky130_fd_sc_hd__dfrtn_1_42/a_639_47# VSS 0.00fF
C17409 sky130_fd_sc_hd__dfrtn_1_42/a_1270_413# VSS 0.00fF
C17410 sky130_fd_sc_hd__dfrtn_1_42/a_651_413# VSS 0.01fF
C17411 sky130_fd_sc_hd__dfrtn_1_42/a_448_47# VSS 0.01fF
C17412 sky130_fd_sc_hd__dfrtn_1_42/a_1108_47# VSS 0.15fF
C17413 sky130_fd_sc_hd__dfrtn_1_42/a_1283_21# VSS 0.29fF
C17414 sky130_fd_sc_hd__dfrtn_1_42/a_543_47# VSS 0.15fF
C17415 sky130_fd_sc_hd__dfrtn_1_42/a_761_289# VSS 0.12fF
C17416 sky130_fd_sc_hd__dfrtn_1_42/a_193_47# VSS 0.26fF
C17417 sky130_fd_sc_hd__dfrtn_1_42/a_27_47# VSS 0.45fF
C17418 sky130_fd_sc_hd__dfrtn_1_31/a_1462_47# VSS 0.00fF
C17419 sky130_fd_sc_hd__dfrtn_1_31/a_1217_47# VSS 0.00fF
C17420 sky130_fd_sc_hd__dfrtn_1_31/a_805_47# VSS 0.00fF
C17421 sky130_fd_sc_hd__dfrtn_1_31/a_639_47# VSS 0.00fF
C17422 sky130_fd_sc_hd__dfrtn_1_31/a_1270_413# VSS 0.00fF
C17423 sky130_fd_sc_hd__dfrtn_1_31/a_651_413# VSS 0.01fF
C17424 sky130_fd_sc_hd__dfrtn_1_31/a_448_47# VSS 0.01fF
C17425 sky130_fd_sc_hd__dfrtn_1_31/a_1108_47# VSS 0.15fF
C17426 sky130_fd_sc_hd__dfrtn_1_31/a_1283_21# VSS 0.29fF
C17427 sky130_fd_sc_hd__dfrtn_1_31/a_543_47# VSS 0.15fF
C17428 sky130_fd_sc_hd__dfrtn_1_31/a_761_289# VSS 0.12fF
C17429 sky130_fd_sc_hd__dfrtn_1_31/a_193_47# VSS 0.14fF
C17430 sky130_fd_sc_hd__dfrtn_1_31/a_27_47# VSS 0.45fF
C17431 sky130_fd_sc_hd__dfrtn_1_20/a_1462_47# VSS 0.00fF
C17432 sky130_fd_sc_hd__dfrtn_1_20/a_1217_47# VSS 0.00fF
C17433 sky130_fd_sc_hd__dfrtn_1_20/a_805_47# VSS 0.00fF
C17434 sky130_fd_sc_hd__dfrtn_1_20/a_639_47# VSS 0.00fF
C17435 sky130_fd_sc_hd__dfrtn_1_20/a_1270_413# VSS 0.00fF
C17436 sky130_fd_sc_hd__dfrtn_1_20/a_651_413# VSS 0.01fF
C17437 sky130_fd_sc_hd__dfrtn_1_20/a_448_47# VSS 0.01fF
C17438 sky130_fd_sc_hd__dfrtn_1_20/a_1108_47# VSS 0.15fF
C17439 sky130_fd_sc_hd__dfrtn_1_20/a_1283_21# VSS 0.29fF
C17440 sky130_fd_sc_hd__dfrtn_1_20/a_543_47# VSS 0.15fF
C17441 sky130_fd_sc_hd__dfrtn_1_20/a_761_289# VSS 0.12fF
C17442 sky130_fd_sc_hd__dfrtn_1_20/a_193_47# VSS 0.24fF
C17443 sky130_fd_sc_hd__dfrtn_1_20/a_27_47# VSS 0.44fF
C17444 sky130_fd_sc_hd__or2_2_0/X VSS 0.13fF
C17445 sky130_fd_sc_hd__dfrtn_1_41/a_1462_47# VSS 0.00fF
C17446 sky130_fd_sc_hd__dfrtn_1_41/a_1217_47# VSS 0.00fF
C17447 sky130_fd_sc_hd__dfrtn_1_41/a_805_47# VSS 0.00fF
C17448 sky130_fd_sc_hd__dfrtn_1_41/a_639_47# VSS 0.00fF
C17449 sky130_fd_sc_hd__dfrtn_1_41/a_1270_413# VSS 0.00fF
C17450 sky130_fd_sc_hd__dfrtn_1_41/a_651_413# VSS 0.01fF
C17451 sky130_fd_sc_hd__dfrtn_1_41/a_448_47# VSS 0.01fF
C17452 sky130_fd_sc_hd__dfrtn_1_41/a_1108_47# VSS 0.15fF
C17453 sky130_fd_sc_hd__dfrtn_1_41/a_1283_21# VSS 0.29fF
C17454 sky130_fd_sc_hd__dfrtn_1_41/a_543_47# VSS 0.15fF
C17455 sky130_fd_sc_hd__dfrtn_1_41/a_761_289# VSS 0.12fF
C17456 sky130_fd_sc_hd__dfrtn_1_41/a_193_47# VSS 0.19fF
C17457 sky130_fd_sc_hd__dfrtn_1_41/a_27_47# VSS 0.41fF
C17458 sky130_fd_sc_hd__dfrtn_1_30/a_1462_47# VSS 0.00fF
C17459 sky130_fd_sc_hd__dfrtn_1_30/a_1217_47# VSS 0.00fF
C17460 sky130_fd_sc_hd__dfrtn_1_30/a_805_47# VSS 0.00fF
C17461 sky130_fd_sc_hd__dfrtn_1_30/a_639_47# VSS 0.00fF
C17462 sky130_fd_sc_hd__dfrtn_1_30/a_1270_413# VSS 0.00fF
C17463 sky130_fd_sc_hd__dfrtn_1_30/a_651_413# VSS 0.01fF
C17464 sky130_fd_sc_hd__dfrtn_1_30/a_448_47# VSS 0.01fF
C17465 sky130_fd_sc_hd__dfrtn_1_30/a_1108_47# VSS 0.15fF
C17466 sky130_fd_sc_hd__dfrtn_1_30/a_1283_21# VSS 0.28fF
C17467 sky130_fd_sc_hd__dfrtn_1_30/a_543_47# VSS 0.15fF
C17468 sky130_fd_sc_hd__dfrtn_1_30/a_761_289# VSS 0.12fF
C17469 sky130_fd_sc_hd__dfrtn_1_30/a_193_47# VSS 0.15fF
C17470 sky130_fd_sc_hd__dfrtn_1_30/a_27_47# VSS 0.43fF
C17471 sky130_fd_sc_hd__dfrtn_1_40/a_1462_47# VSS 0.00fF
C17472 sky130_fd_sc_hd__dfrtn_1_40/a_1217_47# VSS 0.00fF
C17473 sky130_fd_sc_hd__dfrtn_1_40/a_805_47# VSS 0.00fF
C17474 sky130_fd_sc_hd__dfrtn_1_40/a_639_47# VSS 0.00fF
C17475 sky130_fd_sc_hd__dfrtn_1_40/a_1270_413# VSS 0.00fF
C17476 sky130_fd_sc_hd__dfrtn_1_40/a_651_413# VSS 0.00fF
C17477 sky130_fd_sc_hd__dfrtn_1_40/a_448_47# VSS 0.01fF
C17478 sky130_fd_sc_hd__dfrtn_1_40/a_1108_47# VSS 0.15fF
C17479 sky130_fd_sc_hd__dfrtn_1_40/a_1283_21# VSS 0.28fF
C17480 sky130_fd_sc_hd__dfrtn_1_40/a_543_47# VSS 0.15fF
C17481 sky130_fd_sc_hd__dfrtn_1_40/a_761_289# VSS 0.11fF
C17482 sky130_fd_sc_hd__dfrtn_1_40/a_193_47# VSS 0.14fF
C17483 sky130_fd_sc_hd__dfrtn_1_40/a_27_47# VSS 0.42fF
C17484 sky130_fd_sc_hd__inv_1_18/Y VSS 0.15fF
C17485 sky130_fd_sc_hd__nor3_2_1/A VSS 0.37fF
C17486 sky130_fd_sc_hd__o2111a_2_0/a_566_47# VSS 0.05fF
C17487 sky130_fd_sc_hd__o2111a_2_0/a_458_47# VSS 0.00fF
C17488 sky130_fd_sc_hd__o2111a_2_0/a_386_47# VSS 0.00fF
C17489 sky130_fd_sc_hd__o2111a_2_0/a_674_297# VSS 0.00fF
C17490 sky130_fd_sc_hd__o2111a_2_0/a_80_21# VSS 0.27fF
C17491 sky130_fd_sc_hd__nand3b_1_1/a_316_47# VSS 0.00fF
C17492 sky130_fd_sc_hd__nand3b_1_1/a_232_47# VSS 0.00fF
C17493 sky130_fd_sc_hd__nand3b_1_1/a_53_93# VSS 0.23fF
C17494 sky130_fd_sc_hd__or3b_2_0/a_472_297# VSS 0.00fF
C17495 sky130_fd_sc_hd__or3b_2_0/a_388_297# VSS 0.00fF
C17496 sky130_fd_sc_hd__or3b_2_0/a_27_47# VSS 0.23fF
C17497 sky130_fd_sc_hd__or3b_2_0/a_176_21# VSS 0.28fF
C17498 sky130_fd_sc_hd__nor3_2_3/a_281_297# VSS 0.05fF
C17499 sky130_fd_sc_hd__nor3_2_3/a_27_297# VSS 0.07fF
C17500 sky130_fd_sc_hd__nand3b_1_0/a_316_47# VSS 0.00fF
C17501 sky130_fd_sc_hd__nand3b_1_0/a_232_47# VSS 0.00fF
C17502 sky130_fd_sc_hd__nand3b_1_0/a_53_93# VSS 0.22fF
C17503 sky130_fd_sc_hd__nor3_2_2/a_281_297# VSS 0.04fF
C17504 sky130_fd_sc_hd__nor3_2_2/a_27_297# VSS 0.06fF
C17505 sky130_fd_sc_hd__nor3_2_1/a_281_297# VSS 0.05fF
C17506 sky130_fd_sc_hd__nor3_2_1/a_27_297# VSS 0.07fF
C17507 sky130_fd_sc_hd__nor3_2_0/a_281_297# VSS 0.05fF
C17508 sky130_fd_sc_hd__nor3_2_0/a_27_297# VSS 0.07fF
C17509 sky130_fd_sc_hd__nor3_1_19/a_193_297# VSS 0.00fF
C17510 sky130_fd_sc_hd__nor3_1_19/a_109_297# VSS 0.00fF
C17511 sky130_fd_sc_hd__inv_1_54/Y VSS 0.38fF
C17512 sky130_fd_sc_hd__inv_1_33/Y VSS 0.12fF
C17513 sky130_fd_sc_hd__mux4_1_0/a_834_97# VSS 0.03fF
C17514 sky130_fd_sc_hd__mux4_1_0/a_668_97# VSS 0.01fF
C17515 sky130_fd_sc_hd__mux4_1_0/a_193_47# VSS 0.00fF
C17516 sky130_fd_sc_hd__mux4_1_0/a_27_47# VSS 0.07fF
C17517 sky130_fd_sc_hd__mux4_1_0/a_1478_413# VSS 0.17fF
C17518 sky130_fd_sc_hd__mux4_1_0/a_1290_413# VSS 0.24fF
C17519 sky130_fd_sc_hd__mux4_1_0/a_750_97# VSS 0.06fF
C17520 sky130_fd_sc_hd__mux4_1_0/a_757_363# VSS 0.02fF
C17521 sky130_fd_sc_hd__mux4_1_0/a_923_363# VSS 0.00fF
C17522 sky130_fd_sc_hd__mux4_1_0/a_277_47# VSS 0.10fF
C17523 sky130_fd_sc_hd__mux4_1_0/a_247_21# VSS 0.30fF
C17524 sky130_fd_sc_hd__mux4_1_0/a_193_413# VSS 0.01fF
C17525 sky130_fd_sc_hd__mux4_1_0/a_27_413# VSS 0.04fF
C17526 sky130_fd_sc_hd__nor3_1_18/a_193_297# VSS 0.00fF
C17527 sky130_fd_sc_hd__nor3_1_18/a_109_297# VSS 0.00fF
C17528 sky130_fd_sc_hd__inv_1_34/A VSS 0.52fF
C17529 sky130_fd_sc_hd__or2b_1_0/a_301_297# VSS 0.00fF
C17530 sky130_fd_sc_hd__or2b_1_0/a_27_53# VSS 0.17fF
C17531 sky130_fd_sc_hd__or2b_1_0/a_219_297# VSS 0.16fF
C17532 sky130_fd_sc_hd__nor3_1_17/a_193_297# VSS 0.00fF
C17533 sky130_fd_sc_hd__nor3_1_17/a_109_297# VSS 0.00fF
C17534 sky130_fd_sc_hd__nand3b_1_0/Y VSS 0.27fF
C17535 sky130_fd_sc_hd__nor3_1_16/a_193_297# VSS 0.00fF
C17536 sky130_fd_sc_hd__nor3_1_16/a_109_297# VSS 0.00fF
C17537 DOUT[13] VSS 2.81fF
C17538 sky130_fd_sc_hd__inv_1_27/A VSS 0.52fF
C17539 sky130_fd_sc_hd__dfrtp_1_3/a_1462_47# VSS 0.00fF
C17540 sky130_fd_sc_hd__dfrtp_1_3/a_1217_47# VSS 0.00fF
C17541 sky130_fd_sc_hd__dfrtp_1_3/a_805_47# VSS 0.00fF
C17542 sky130_fd_sc_hd__dfrtp_1_3/a_639_47# VSS 0.00fF
C17543 sky130_fd_sc_hd__dfrtp_1_3/a_1270_413# VSS 0.00fF
C17544 sky130_fd_sc_hd__dfrtp_1_3/a_651_413# VSS 0.01fF
C17545 sky130_fd_sc_hd__dfrtp_1_3/a_448_47# VSS 0.02fF
C17546 sky130_fd_sc_hd__dfrtp_1_3/a_1108_47# VSS 0.16fF
C17547 sky130_fd_sc_hd__dfrtp_1_3/a_1283_21# VSS 0.30fF
C17548 sky130_fd_sc_hd__dfrtp_1_3/a_543_47# VSS 0.16fF
C17549 sky130_fd_sc_hd__dfrtp_1_3/a_761_289# VSS 0.13fF
C17550 sky130_fd_sc_hd__dfrtp_1_3/a_193_47# VSS 0.28fF
C17551 sky130_fd_sc_hd__dfrtp_1_3/a_27_47# VSS 0.33fF
C17552 sky130_fd_sc_hd__nor3_1_15/a_193_297# VSS 0.00fF
C17553 sky130_fd_sc_hd__nor3_1_15/a_109_297# VSS 0.00fF
C17554 CLK_REF VSS 2.38fF
C17555 sky130_fd_sc_hd__dfrtp_1_2/a_1462_47# VSS 0.00fF
C17556 sky130_fd_sc_hd__dfrtp_1_2/a_1217_47# VSS 0.00fF
C17557 sky130_fd_sc_hd__dfrtp_1_2/a_805_47# VSS 0.00fF
C17558 sky130_fd_sc_hd__dfrtp_1_2/a_639_47# VSS 0.00fF
C17559 sky130_fd_sc_hd__dfrtp_1_2/a_1270_413# VSS 0.00fF
C17560 sky130_fd_sc_hd__dfrtp_1_2/a_651_413# VSS 0.01fF
C17561 sky130_fd_sc_hd__dfrtp_1_2/a_448_47# VSS 0.02fF
C17562 sky130_fd_sc_hd__dfrtp_1_2/a_1108_47# VSS 0.15fF
C17563 sky130_fd_sc_hd__dfrtp_1_2/a_1283_21# VSS 0.29fF
C17564 sky130_fd_sc_hd__dfrtp_1_2/a_543_47# VSS 0.15fF
C17565 sky130_fd_sc_hd__dfrtp_1_2/a_761_289# VSS 0.12fF
C17566 sky130_fd_sc_hd__dfrtp_1_2/a_193_47# VSS 0.27fF
C17567 sky130_fd_sc_hd__dfrtp_1_2/a_27_47# VSS 0.30fF
C17568 sky130_fd_sc_hd__nor3_1_14/a_193_297# VSS 0.00fF
C17569 sky130_fd_sc_hd__nor3_1_14/a_109_297# VSS 0.00fF
C17570 sky130_fd_sc_hd__inv_1_30/A VSS 0.66fF
C17571 sky130_fd_sc_hd__nor2_1_0/a_109_297# VSS -0.00fF
C17572 sky130_fd_sc_hd__dfrtp_1_1/a_1462_47# VSS 0.00fF
C17573 sky130_fd_sc_hd__dfrtp_1_1/a_1217_47# VSS 0.00fF
C17574 sky130_fd_sc_hd__dfrtp_1_1/a_805_47# VSS 0.00fF
C17575 sky130_fd_sc_hd__dfrtp_1_1/a_639_47# VSS 0.00fF
C17576 sky130_fd_sc_hd__dfrtp_1_1/a_1270_413# VSS 0.00fF
C17577 sky130_fd_sc_hd__dfrtp_1_1/a_651_413# VSS 0.01fF
C17578 sky130_fd_sc_hd__dfrtp_1_1/a_448_47# VSS 0.02fF
C17579 sky130_fd_sc_hd__dfrtp_1_1/a_1108_47# VSS 0.17fF
C17580 sky130_fd_sc_hd__dfrtp_1_1/a_1283_21# VSS 0.31fF
C17581 sky130_fd_sc_hd__dfrtp_1_1/a_543_47# VSS 0.16fF
C17582 sky130_fd_sc_hd__dfrtp_1_1/a_761_289# VSS 0.13fF
C17583 sky130_fd_sc_hd__dfrtp_1_1/a_193_47# VSS 0.30fF
C17584 sky130_fd_sc_hd__dfrtp_1_1/a_27_47# VSS 0.45fF
C17585 sky130_fd_sc_hd__nor3_1_13/a_193_297# VSS 0.00fF
C17586 sky130_fd_sc_hd__nor3_1_13/a_109_297# VSS 0.00fF
C17587 sky130_fd_sc_hd__inv_1_29/A VSS 2.19fF
C17588 sky130_fd_sc_hd__a221oi_4_0/a_1241_47# VSS 0.02fF
C17589 sky130_fd_sc_hd__a221oi_4_0/a_453_47# VSS 0.01fF
C17590 sky130_fd_sc_hd__a221oi_4_0/a_471_297# VSS 0.07fF
C17591 sky130_fd_sc_hd__a221oi_4_0/a_27_297# VSS 0.07fF
C17592 sky130_fd_sc_hd__dfrtp_1_0/a_1462_47# VSS 0.00fF
C17593 sky130_fd_sc_hd__dfrtp_1_0/a_1217_47# VSS 0.00fF
C17594 sky130_fd_sc_hd__dfrtp_1_0/a_805_47# VSS 0.00fF
C17595 sky130_fd_sc_hd__dfrtp_1_0/a_639_47# VSS 0.00fF
C17596 sky130_fd_sc_hd__dfrtp_1_0/a_1270_413# VSS 0.00fF
C17597 sky130_fd_sc_hd__dfrtp_1_0/a_651_413# VSS 0.01fF
C17598 sky130_fd_sc_hd__dfrtp_1_0/a_448_47# VSS 0.02fF
C17599 sky130_fd_sc_hd__dfrtp_1_0/a_1108_47# VSS 0.16fF
C17600 sky130_fd_sc_hd__dfrtp_1_0/a_1283_21# VSS 0.30fF
C17601 sky130_fd_sc_hd__dfrtp_1_0/a_543_47# VSS 0.16fF
C17602 sky130_fd_sc_hd__dfrtp_1_0/a_761_289# VSS 0.12fF
C17603 sky130_fd_sc_hd__dfrtp_1_0/a_193_47# VSS 0.28fF
C17604 sky130_fd_sc_hd__dfrtp_1_0/a_27_47# VSS 0.46fF
C17605 sky130_fd_sc_hd__inv_1_4/A VSS 0.36fF
C17606 sky130_fd_sc_hd__nor3_1_12/a_193_297# VSS 0.00fF
C17607 sky130_fd_sc_hd__nor3_1_12/a_109_297# VSS 0.00fF
C17608 sky130_fd_sc_hd__inv_1_52/A VSS 2.61fF
C17609 sky130_fd_sc_hd__nor3_1_9/a_193_297# VSS 0.00fF
C17610 sky130_fd_sc_hd__nor3_1_9/a_109_297# VSS 0.00fF
C17611 sky130_fd_sc_hd__inv_1_10/A VSS 1.25fF
C17612 sky130_fd_sc_hd__nor3_1_11/a_193_297# VSS 0.00fF
C17613 sky130_fd_sc_hd__nor3_1_11/a_109_297# VSS 0.00fF
C17614 sky130_fd_sc_hd__inv_1_49/Y VSS 0.12fF
C17615 sky130_fd_sc_hd__nor3_1_8/a_193_297# VSS 0.00fF
C17616 sky130_fd_sc_hd__nor3_1_8/a_109_297# VSS 0.00fF
C17617 sky130_fd_sc_hd__nor3_1_10/a_193_297# VSS 0.00fF
C17618 sky130_fd_sc_hd__nor3_1_10/a_109_297# VSS 0.00fF
C17619 sky130_fd_sc_hd__nor3_1_7/a_193_297# VSS 0.00fF
C17620 sky130_fd_sc_hd__nor3_1_7/a_109_297# VSS 0.00fF
C17621 sky130_fd_sc_hd__inv_1_0/A VSS 0.37fF
C17622 HEADER_2/a_508_138# VSS 0.16fF
C17623 sky130_fd_sc_hd__nor3_1_20/a_193_297# VSS 0.00fF
C17624 sky130_fd_sc_hd__nor3_1_20/a_109_297# VSS 0.00fF
C17625 sky130_fd_sc_hd__mux4_2_0/X VSS 0.22fF
C17626 sky130_fd_sc_hd__nor3_1_6/a_193_297# VSS 0.00fF
C17627 sky130_fd_sc_hd__nor3_1_6/a_109_297# VSS 0.00fF
C17628 sky130_fd_sc_hd__or3_1_0/a_183_297# VSS 0.00fF
C17629 sky130_fd_sc_hd__or3_1_0/a_111_297# VSS 0.00fF
C17630 sky130_fd_sc_hd__or3_1_0/a_29_53# VSS 0.21fF
C17631 HEADER_1/a_508_138# VSS 0.16fF
.ends

